module SRAMTemplate(
  input         clock,
  input         reset,
  output        io_r_req_ready,
  input         io_r_req_valid,
  input  [8:0]  io_r_req_bits_setIdx,
  output [27:0] io_r_resp_data_0_tag,
  output [1:0]  io_r_resp_data_0__type,
  output [38:0] io_r_resp_data_0_target,
  output [2:0]  io_r_resp_data_0_brIdx,
  output        io_r_resp_data_0_valid,
  input         io_w_req_valid,
  input  [8:0]  io_w_req_bits_setIdx,
  input  [27:0] io_w_req_bits_data_tag,
  input  [1:0]  io_w_req_bits_data__type,
  input  [38:0] io_w_req_bits_data_target,
  input  [2:0]  io_w_req_bits_data_brIdx
);
`ifdef RANDOMIZE_MEM_INIT
  reg [95:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [95:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [72:0] array_0 [0:511]; // @[SRAMTemplate.scala 76:26]
  wire [72:0] array_0__T_19_data; // @[SRAMTemplate.scala 76:26]
  wire [8:0] array_0__T_19_addr; // @[SRAMTemplate.scala 76:26]
  wire [72:0] array_0__T_15_data; // @[SRAMTemplate.scala 76:26]
  wire [8:0] array_0__T_15_addr; // @[SRAMTemplate.scala 76:26]
  wire  array_0__T_15_mask; // @[SRAMTemplate.scala 76:26]
  wire  array_0__T_15_en; // @[SRAMTemplate.scala 76:26]
  reg  array_0__T_19_en_pipe_0;
  reg [8:0] array_0__T_19_addr_pipe_0;
  reg  resetState; // @[SRAMTemplate.scala 80:30]
  reg [8:0] resetSet; // @[Counter.scala 29:33]
  wire  _T_3 = resetSet == 9'h1ff; // @[Counter.scala 38:24]
  wire [8:0] _T_5 = resetSet + 9'h1; // @[Counter.scala 39:22]
  wire  _GEN_1 = resetState & _T_3; // @[Counter.scala 67:17]
  wire  _GEN_2 = _GEN_1 ? 1'h0 : resetState; // @[SRAMTemplate.scala 82:24]
  wire  wen = io_w_req_valid | resetState; // @[SRAMTemplate.scala 88:52]
  wire  _T_6 = ~wen; // @[SRAMTemplate.scala 89:41]
  wire [72:0] _T_11 = {io_w_req_bits_data_tag,io_w_req_bits_data__type,io_w_req_bits_data_target,io_w_req_bits_data_brIdx,1'h1}; // @[SRAMTemplate.scala 92:78]
  reg  _T_20; // @[Hold.scala 28:106]
  reg [72:0] _T_22_0; // @[Reg.scala 27:20]
  wire [72:0] _GEN_14 = _T_20 ? array_0__T_19_data : _T_22_0; // @[Reg.scala 28:19]
  wire  _T_31 = ~resetState; // @[SRAMTemplate.scala 101:21]
  assign array_0__T_19_addr = array_0__T_19_addr_pipe_0;
  assign array_0__T_19_data = array_0[array_0__T_19_addr]; // @[SRAMTemplate.scala 76:26]
  assign array_0__T_15_data = resetState ? 73'h0 : _T_11;
  assign array_0__T_15_addr = resetState ? resetSet : io_w_req_bits_setIdx;
  assign array_0__T_15_mask = 1'h1;
  assign array_0__T_15_en = io_w_req_valid | resetState;
  assign io_r_req_ready = _T_31 & _T_6; // @[SRAMTemplate.scala 101:18]
  assign io_r_resp_data_0_tag = _GEN_14[72:45]; // @[SRAMTemplate.scala 99:18]
  assign io_r_resp_data_0__type = _GEN_14[44:43]; // @[SRAMTemplate.scala 99:18]
  assign io_r_resp_data_0_target = _GEN_14[42:4]; // @[SRAMTemplate.scala 99:18]
  assign io_r_resp_data_0_brIdx = _GEN_14[3:1]; // @[SRAMTemplate.scala 99:18]
  assign io_r_resp_data_0_valid = _GEN_14[0]; // @[SRAMTemplate.scala 99:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {3{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    array_0[initvar] = _RAND_0[72:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  array_0__T_19_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  array_0__T_19_addr_pipe_0 = _RAND_2[8:0];
  _RAND_3 = {1{`RANDOM}};
  resetState = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  resetSet = _RAND_4[8:0];
  _RAND_5 = {1{`RANDOM}};
  _T_20 = _RAND_5[0:0];
  _RAND_6 = {3{`RANDOM}};
  _T_22_0 = _RAND_6[72:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(array_0__T_15_en & array_0__T_15_mask) begin
      array_0[array_0__T_15_addr] <= array_0__T_15_data; // @[SRAMTemplate.scala 76:26]
    end
    array_0__T_19_en_pipe_0 <= io_r_req_valid & _T_6;
    if (io_r_req_valid & _T_6) begin
      array_0__T_19_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    resetState <= reset | _GEN_2;
    if (reset) begin
      resetSet <= 9'h0;
    end else if (resetState) begin
      resetSet <= _T_5;
    end
    _T_20 <= io_r_req_valid & _T_6;
    if (reset) begin
      _T_22_0 <= 73'h0;
    end else if (_T_20) begin
      _T_22_0 <= array_0__T_19_data;
    end
  end
endmodule
module BPU_inorder(
  input         clock,
  input         reset,
  input         io_in_pc_valid,
  input  [38:0] io_in_pc_bits,
  output [38:0] io_out_target,
  output        io_out_valid,
  input         io_flush,
  output [2:0]  io_brIdx,
  output        io_crosslineJump,
  input         MOUFlushICache,
  input         bpuUpdateReq_valid,
  input  [38:0] bpuUpdateReq_pc,
  input         bpuUpdateReq_isMissPredict,
  input  [38:0] bpuUpdateReq_actualTarget,
  input         bpuUpdateReq_actualTaken,
  input  [6:0]  bpuUpdateReq_fuOpType,
  input  [1:0]  bpuUpdateReq_btbType,
  input         bpuUpdateReq_isRVC,
  input         DISPLAY_ENABLE,
  input         MOUFlushTLB
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire  btb_clock; // @[BPU.scala 302:19]
  wire  btb_reset; // @[BPU.scala 302:19]
  wire  btb_io_r_req_ready; // @[BPU.scala 302:19]
  wire  btb_io_r_req_valid; // @[BPU.scala 302:19]
  wire [8:0] btb_io_r_req_bits_setIdx; // @[BPU.scala 302:19]
  wire [27:0] btb_io_r_resp_data_0_tag; // @[BPU.scala 302:19]
  wire [1:0] btb_io_r_resp_data_0__type; // @[BPU.scala 302:19]
  wire [38:0] btb_io_r_resp_data_0_target; // @[BPU.scala 302:19]
  wire [2:0] btb_io_r_resp_data_0_brIdx; // @[BPU.scala 302:19]
  wire  btb_io_r_resp_data_0_valid; // @[BPU.scala 302:19]
  wire  btb_io_w_req_valid; // @[BPU.scala 302:19]
  wire [8:0] btb_io_w_req_bits_setIdx; // @[BPU.scala 302:19]
  wire [27:0] btb_io_w_req_bits_data_tag; // @[BPU.scala 302:19]
  wire [1:0] btb_io_w_req_bits_data__type; // @[BPU.scala 302:19]
  wire [38:0] btb_io_w_req_bits_data_target; // @[BPU.scala 302:19]
  wire [2:0] btb_io_w_req_bits_data_brIdx; // @[BPU.scala 302:19]
  reg [1:0] pht [0:511]; // @[BPU.scala 336:16]
  wire [1:0] pht__T_81_data; // @[BPU.scala 336:16]
  wire [8:0] pht__T_81_addr; // @[BPU.scala 336:16]
  wire [1:0] pht__T_139_data; // @[BPU.scala 336:16]
  wire [8:0] pht__T_139_addr; // @[BPU.scala 336:16]
  wire [1:0] pht__T_160_data; // @[BPU.scala 336:16]
  wire [8:0] pht__T_160_addr; // @[BPU.scala 336:16]
  wire  pht__T_160_mask; // @[BPU.scala 336:16]
  wire  pht__T_160_en; // @[BPU.scala 336:16]
  reg [38:0] ras [0:15]; // @[BPU.scala 342:16]
  wire [38:0] ras__T_83_data; // @[BPU.scala 342:16]
  wire [3:0] ras__T_83_addr; // @[BPU.scala 342:16]
  wire [38:0] ras__T_169_data; // @[BPU.scala 342:16]
  wire [3:0] ras__T_169_addr; // @[BPU.scala 342:16]
  wire  ras__T_169_mask; // @[BPU.scala 342:16]
  wire  ras__T_169_en; // @[BPU.scala 342:16]
  reg  flush; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = io_in_pc_valid ? 1'h0 : flush; // @[StopWatch.scala 26:19]
  wire  _GEN_1 = io_flush | _GEN_0; // @[StopWatch.scala 27:20]
  wire  _T_1 = MOUFlushICache | MOUFlushTLB; // @[BPU.scala 308:42]
  wire  _T_2 = reset | _T_1; // @[BPU.scala 308:29]
  reg [63:0] _T_6; // @[GTimer.scala 24:20]
  wire [63:0] _T_8 = _T_6 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_10 = _T_2 & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  wire  _T_12 = ~reset; // @[Debug.scala 56:24]
  reg [38:0] pcLatch; // @[Reg.scala 15:16]
  wire [27:0] btbRead_tag = btb_io_r_resp_data_0_tag; // @[BPU.scala 315:21 BPU.scala 316:11]
  wire  _T_27 = btbRead_tag == pcLatch[38:11]; // @[BPU.scala 320:45]
  wire  btbRead_valid = btb_io_r_resp_data_0_valid; // @[BPU.scala 315:21 BPU.scala 316:11]
  wire  _T_28 = btbRead_valid & _T_27; // @[BPU.scala 320:30]
  wire  _T_29 = ~flush; // @[BPU.scala 320:76]
  wire  _T_30 = _T_28 & _T_29; // @[BPU.scala 320:73]
  wire  _T_31 = btb_io_r_req_ready & btb_io_r_req_valid; // @[Decoupled.scala 40:37]
  reg  _T_32; // @[BPU.scala 320:93]
  wire  _T_33 = _T_30 & _T_32; // @[BPU.scala 320:83]
  wire [2:0] btbRead_brIdx = btb_io_r_resp_data_0_brIdx; // @[BPU.scala 315:21 BPU.scala 316:11]
  wire  _T_36 = pcLatch[1] & btbRead_brIdx[0]; // @[BPU.scala 320:147]
  wire  _T_37 = ~_T_36; // @[BPU.scala 320:134]
  wire  btbHit = _T_33 & _T_37; // @[BPU.scala 320:131]
  wire  crosslineJump = btbRead_brIdx[2] & btbHit; // @[BPU.scala 327:40]
  reg [63:0] _T_39; // @[GTimer.scala 24:20]
  wire [63:0] _T_41 = _T_39 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_54; // @[GTimer.scala 24:20]
  wire [63:0] _T_56 = _T_54 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_58 = btbHit & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  wire [1:0] _T_64 = io_out_valid ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [2:0] _T_65 = {crosslineJump,_T_64}; // @[Cat.scala 29:58]
  reg [63:0] _T_66; // @[GTimer.scala 24:20]
  wire [63:0] _T_68 = _T_66 + 64'h1; // @[GTimer.scala 25:12]
  reg  phtTaken; // @[Reg.scala 15:16]
  reg [3:0] value; // @[Counter.scala 29:33]
  reg [38:0] rasTarget; // @[Reg.scala 15:16]
  wire  _T_100 = ~bpuUpdateReq_pc[1]; // @[BPU.scala 353:150]
  wire [1:0] _T_101 = {bpuUpdateReq_pc[1],_T_100}; // @[Cat.scala 29:58]
  reg [63:0] _T_102; // @[GTimer.scala 24:20]
  wire [63:0] _T_104 = _T_102 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_106 = bpuUpdateReq_valid & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  wire  _T_118 = bpuUpdateReq_pc[2:0] == 3'h6; // @[BPU.scala 367:36]
  wire  _T_119 = ~bpuUpdateReq_isRVC; // @[BPU.scala 367:49]
  wire  _T_120 = _T_118 & _T_119; // @[BPU.scala 367:46]
  wire [1:0] _T_124 = {_T_120,bpuUpdateReq_pc[1]}; // @[Cat.scala 29:58]
  reg [1:0] cnt; // @[BPU.scala 389:20]
  reg  reqLatch_valid; // @[BPU.scala 390:25]
  reg [38:0] reqLatch_pc; // @[BPU.scala 390:25]
  reg  reqLatch_actualTaken; // @[BPU.scala 390:25]
  reg [6:0] reqLatch_fuOpType; // @[BPU.scala 390:25]
  wire  _T_141 = ~reqLatch_fuOpType[3]; // @[ALU.scala 62:30]
  wire  _T_142 = reqLatch_valid & _T_141; // @[BPU.scala 391:24]
  wire [1:0] _T_144 = cnt + 2'h1; // @[BPU.scala 393:33]
  wire [1:0] _T_146 = cnt - 2'h1; // @[BPU.scala 393:44]
  wire  _T_148 = cnt != 2'h3; // @[BPU.scala 394:30]
  wire  _T_149 = reqLatch_actualTaken & _T_148; // @[BPU.scala 394:22]
  wire  _T_150 = ~reqLatch_actualTaken; // @[BPU.scala 394:48]
  wire  _T_151 = cnt != 2'h0; // @[BPU.scala 394:63]
  wire  _T_152 = _T_150 & _T_151; // @[BPU.scala 394:55]
  wire  _T_153 = _T_149 | _T_152; // @[BPU.scala 394:44]
  wire  _T_161 = bpuUpdateReq_fuOpType == 7'h5c; // @[BPU.scala 403:24]
  wire [3:0] _T_163 = value + 4'h1; // @[BPU.scala 404:26]
  wire [38:0] _T_165 = bpuUpdateReq_pc + 39'h2; // @[BPU.scala 404:55]
  wire [38:0] _T_167 = bpuUpdateReq_pc + 39'h4; // @[BPU.scala 404:69]
  wire  _T_172 = bpuUpdateReq_fuOpType == 7'h5e; // @[BPU.scala 408:29]
  wire  _T_173 = value == 4'h0; // @[BPU.scala 409:21]
  wire [3:0] _T_176 = value - 4'h1; // @[BPU.scala 412:53]
  wire [1:0] btbRead__type = btb_io_r_resp_data_0__type; // @[BPU.scala 315:21 BPU.scala 316:11]
  wire  _T_178 = btbRead__type == 2'h3; // @[BPU.scala 416:38]
  wire [38:0] btbRead_target = btb_io_r_resp_data_0_target; // @[BPU.scala 315:21 BPU.scala 316:11]
  wire [3:0] _T_183 = {1'h1,crosslineJump,_T_64}; // @[Cat.scala 29:58]
  wire [3:0] _GEN_28 = {{1'd0}, btbRead_brIdx}; // @[BPU.scala 419:30]
  wire [3:0] _T_184 = _GEN_28 & _T_183; // @[BPU.scala 419:30]
  wire  _T_185 = btbRead__type == 2'h0; // @[BPU.scala 420:47]
  wire  _T_186 = rasTarget != 39'h0; // @[BPU.scala 420:91]
  wire  _T_188 = _T_185 ? phtTaken : _T_186; // @[BPU.scala 420:32]
  SRAMTemplate btb ( // @[BPU.scala 302:19]
    .clock(btb_clock),
    .reset(btb_reset),
    .io_r_req_ready(btb_io_r_req_ready),
    .io_r_req_valid(btb_io_r_req_valid),
    .io_r_req_bits_setIdx(btb_io_r_req_bits_setIdx),
    .io_r_resp_data_0_tag(btb_io_r_resp_data_0_tag),
    .io_r_resp_data_0__type(btb_io_r_resp_data_0__type),
    .io_r_resp_data_0_target(btb_io_r_resp_data_0_target),
    .io_r_resp_data_0_brIdx(btb_io_r_resp_data_0_brIdx),
    .io_r_resp_data_0_valid(btb_io_r_resp_data_0_valid),
    .io_w_req_valid(btb_io_w_req_valid),
    .io_w_req_bits_setIdx(btb_io_w_req_bits_setIdx),
    .io_w_req_bits_data_tag(btb_io_w_req_bits_data_tag),
    .io_w_req_bits_data__type(btb_io_w_req_bits_data__type),
    .io_w_req_bits_data_target(btb_io_w_req_bits_data_target),
    .io_w_req_bits_data_brIdx(btb_io_w_req_bits_data_brIdx)
  );
  assign pht__T_81_addr = io_in_pc_bits[10:2];
  assign pht__T_81_data = pht[pht__T_81_addr]; // @[BPU.scala 336:16]
  assign pht__T_139_addr = bpuUpdateReq_pc[10:2];
  assign pht__T_139_data = pht[pht__T_139_addr]; // @[BPU.scala 336:16]
  assign pht__T_160_data = reqLatch_actualTaken ? _T_144 : _T_146;
  assign pht__T_160_addr = reqLatch_pc[10:2];
  assign pht__T_160_mask = 1'h1;
  assign pht__T_160_en = _T_142 & _T_153;
  assign ras__T_83_addr = value;
  assign ras__T_83_data = ras[ras__T_83_addr]; // @[BPU.scala 342:16]
  assign ras__T_169_data = bpuUpdateReq_isRVC ? _T_165 : _T_167;
  assign ras__T_169_addr = value + 4'h1;
  assign ras__T_169_mask = 1'h1;
  assign ras__T_169_en = bpuUpdateReq_valid & _T_161;
  assign io_out_target = _T_178 ? rasTarget : btbRead_target; // @[BPU.scala 416:17]
  assign io_out_valid = btbHit & _T_188; // @[BPU.scala 420:16]
  assign io_brIdx = _T_184[2:0]; // @[BPU.scala 419:13]
  assign io_crosslineJump = btbRead_brIdx[2] & btbHit; // @[BPU.scala 328:20]
  assign btb_clock = clock;
  assign btb_reset = reset | _T_1; // @[BPU.scala 308:13]
  assign btb_io_r_req_valid = io_in_pc_valid; // @[BPU.scala 311:22]
  assign btb_io_r_req_bits_setIdx = io_in_pc_bits[10:2]; // @[BPU.scala 312:28]
  assign btb_io_w_req_valid = bpuUpdateReq_isMissPredict & bpuUpdateReq_valid; // @[BPU.scala 375:22]
  assign btb_io_w_req_bits_setIdx = bpuUpdateReq_pc[10:2]; // @[BPU.scala 376:28]
  assign btb_io_w_req_bits_data_tag = bpuUpdateReq_pc[38:11]; // @[BPU.scala 377:26]
  assign btb_io_w_req_bits_data__type = bpuUpdateReq_btbType; // @[BPU.scala 377:26]
  assign btb_io_w_req_bits_data_target = bpuUpdateReq_actualTarget; // @[BPU.scala 377:26]
  assign btb_io_w_req_bits_data_brIdx = {_T_124,_T_100}; // @[BPU.scala 377:26]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    pht[initvar] = _RAND_0[1:0];
  _RAND_1 = {2{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ras[initvar] = _RAND_1[38:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  flush = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  _T_6 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  pcLatch = _RAND_4[38:0];
  _RAND_5 = {1{`RANDOM}};
  _T_32 = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  _T_39 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  _T_54 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  _T_66 = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  phtTaken = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  value = _RAND_10[3:0];
  _RAND_11 = {2{`RANDOM}};
  rasTarget = _RAND_11[38:0];
  _RAND_12 = {2{`RANDOM}};
  _T_102 = _RAND_12[63:0];
  _RAND_13 = {1{`RANDOM}};
  cnt = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  reqLatch_valid = _RAND_14[0:0];
  _RAND_15 = {2{`RANDOM}};
  reqLatch_pc = _RAND_15[38:0];
  _RAND_16 = {1{`RANDOM}};
  reqLatch_actualTaken = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  reqLatch_fuOpType = _RAND_17[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(pht__T_160_en & pht__T_160_mask) begin
      pht[pht__T_160_addr] <= pht__T_160_data; // @[BPU.scala 336:16]
    end
    if(ras__T_169_en & ras__T_169_mask) begin
      ras[ras__T_169_addr] <= ras__T_169_data; // @[BPU.scala 342:16]
    end
    if (reset) begin
      flush <= 1'h0;
    end else begin
      flush <= _GEN_1;
    end
    if (reset) begin
      _T_6 <= 64'h0;
    end else begin
      _T_6 <= _T_8;
    end
    if (io_in_pc_valid) begin
      pcLatch <= io_in_pc_bits;
    end
    if (reset) begin
      _T_32 <= 1'h0;
    end else begin
      _T_32 <= _T_31;
    end
    if (reset) begin
      _T_39 <= 64'h0;
    end else begin
      _T_39 <= _T_41;
    end
    if (reset) begin
      _T_54 <= 64'h0;
    end else begin
      _T_54 <= _T_56;
    end
    if (reset) begin
      _T_66 <= 64'h0;
    end else begin
      _T_66 <= _T_68;
    end
    if (io_in_pc_valid) begin
      phtTaken <= pht__T_81_data[1];
    end
    if (reset) begin
      value <= 4'h0;
    end else if (bpuUpdateReq_valid) begin
      if (_T_161) begin
        value <= _T_163;
      end else if (_T_172) begin
        if (_T_173) begin
          value <= 4'h0;
        end else begin
          value <= _T_176;
        end
      end
    end
    if (io_in_pc_valid) begin
      rasTarget <= ras__T_83_data;
    end
    if (reset) begin
      _T_102 <= 64'h0;
    end else begin
      _T_102 <= _T_104;
    end
    cnt <= pht__T_139_data;
    reqLatch_valid <= bpuUpdateReq_valid;
    reqLatch_pc <= bpuUpdateReq_pc;
    reqLatch_actualTaken <= bpuUpdateReq_actualTaken;
    reqLatch_fuOpType <= bpuUpdateReq_fuOpType;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & _T_12) begin
          $fwrite(32'h80000002,"[%d] BPU_inorder: ",_T_6); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & _T_12) begin
          $fwrite(32'h80000002,"[BPU-RESET] bpu-reset flushBTB:%d flushTLB:%d\n",MOUFlushICache,MOUFlushTLB); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_58 & _T_12) begin
          $fwrite(32'h80000002,"[%d] BPU_inorder: ",_T_54); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_58 & _T_12) begin
          $fwrite(32'h80000002,"[BTBHT1] %d pc=%x tag=%x,%x index=%x bridx=%x tgt=%x,%x flush %x type:%x\n",_T_39,pcLatch,btbRead_tag,pcLatch[38:11],pcLatch[10:2],btbRead_brIdx,btbRead_target,io_out_target,flush,btbRead__type); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_58 & _T_12) begin
          $fwrite(32'h80000002,"[%d] BPU_inorder: ",_T_66); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_58 & _T_12) begin
          $fwrite(32'h80000002,"[BTBHT2] btbRead.brIdx %x mask %x\n",btbRead_brIdx,_T_65); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_106 & _T_12) begin
          $fwrite(32'h80000002,"[%d] BPU_inorder: ",_T_102); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_106 & _T_12) begin
          $fwrite(32'h80000002,"[BTBUP] pc=%x tag=%x index=%x bridx=%x tgt=%x type=%x\n",bpuUpdateReq_pc,bpuUpdateReq_pc[38:11],bpuUpdateReq_pc[10:2],_T_101,bpuUpdateReq_actualTarget,bpuUpdateReq_btbType); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module IFU_inorder(
  input         clock,
  input         reset,
  input         io_imem_req_ready,
  output        io_imem_req_valid,
  output [38:0] io_imem_req_bits_addr,
  output [81:0] io_imem_req_bits_user,
  output        io_imem_resp_ready,
  input         io_imem_resp_valid,
  input  [63:0] io_imem_resp_bits_rdata,
  input  [81:0] io_imem_resp_bits_user,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_instr,
  output [38:0] io_out_bits_pc,
  output [38:0] io_out_bits_pnpc,
  output        io_out_bits_exceptionVec_12,
  output [3:0]  io_out_bits_brIdx,
  input  [38:0] io_redirect_target,
  input         io_redirect_valid,
  output [3:0]  io_flushVec,
  input         io_ipf,
  input         flushICache,
  input         _T_243_valid,
  input  [38:0] _T_243_pc,
  input         _T_243_isMissPredict,
  input  [38:0] _T_243_actualTarget,
  input         _T_243_actualTaken,
  input  [6:0]  _T_243_fuOpType,
  input  [1:0]  _T_243_btbType,
  input         _T_243_isRVC,
  input         DISPLAY_ENABLE,
  output        _T_65_0,
  input         flushTLB,
  output        _T_66_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  bp1_clock; // @[IFU.scala 325:19]
  wire  bp1_reset; // @[IFU.scala 325:19]
  wire  bp1_io_in_pc_valid; // @[IFU.scala 325:19]
  wire [38:0] bp1_io_in_pc_bits; // @[IFU.scala 325:19]
  wire [38:0] bp1_io_out_target; // @[IFU.scala 325:19]
  wire  bp1_io_out_valid; // @[IFU.scala 325:19]
  wire  bp1_io_flush; // @[IFU.scala 325:19]
  wire [2:0] bp1_io_brIdx; // @[IFU.scala 325:19]
  wire  bp1_io_crosslineJump; // @[IFU.scala 325:19]
  wire  bp1_MOUFlushICache; // @[IFU.scala 325:19]
  wire  bp1_bpuUpdateReq_valid; // @[IFU.scala 325:19]
  wire [38:0] bp1_bpuUpdateReq_pc; // @[IFU.scala 325:19]
  wire  bp1_bpuUpdateReq_isMissPredict; // @[IFU.scala 325:19]
  wire [38:0] bp1_bpuUpdateReq_actualTarget; // @[IFU.scala 325:19]
  wire  bp1_bpuUpdateReq_actualTaken; // @[IFU.scala 325:19]
  wire [6:0] bp1_bpuUpdateReq_fuOpType; // @[IFU.scala 325:19]
  wire [1:0] bp1_bpuUpdateReq_btbType; // @[IFU.scala 325:19]
  wire  bp1_bpuUpdateReq_isRVC; // @[IFU.scala 325:19]
  wire  bp1_DISPLAY_ENABLE; // @[IFU.scala 325:19]
  wire  bp1_MOUFlushTLB; // @[IFU.scala 325:19]
  reg [38:0] pc; // @[IFU.scala 321:19]
  wire  _T = io_imem_req_ready & io_imem_req_valid; // @[Decoupled.scala 40:37]
  wire  pcUpdate = io_redirect_valid | _T; // @[IFU.scala 322:36]
  wire [38:0] _T_3 = pc + 39'h2; // @[IFU.scala 323:28]
  wire [38:0] _T_5 = pc + 39'h4; // @[IFU.scala 323:38]
  wire [38:0] snpc = pc[1] ? _T_3 : _T_5; // @[IFU.scala 323:17]
  reg  crosslineJumpLatch; // @[IFU.scala 328:35]
  wire  _T_6 = pcUpdate | bp1_io_flush; // @[IFU.scala 329:17]
  wire  _T_7 = ~crosslineJumpLatch; // @[IFU.scala 330:71]
  wire  _T_8 = bp1_io_crosslineJump & _T_7; // @[IFU.scala 330:68]
  reg [38:0] crosslineJumpTarget; // @[Reg.scala 15:16]
  wire [38:0] pnpc = bp1_io_crosslineJump ? snpc : bp1_io_out_target; // @[IFU.scala 337:17]
  wire [38:0] _T_11 = bp1_io_out_valid ? pnpc : snpc; // @[IFU.scala 339:104]
  wire [38:0] _T_12 = crosslineJumpLatch ? crosslineJumpTarget : _T_11; // @[IFU.scala 339:59]
  wire [38:0] npc = io_redirect_valid ? io_redirect_target : _T_12; // @[IFU.scala 339:16]
  wire  _T_13 = bp1_io_out_valid ? 1'h0 : 1'h1; // @[IFU.scala 340:114]
  wire  _T_14 = bp1_io_crosslineJump | _T_13; // @[IFU.scala 340:87]
  wire  _T_15 = crosslineJumpLatch ? 1'h0 : _T_14; // @[IFU.scala 340:54]
  wire  npcIsSeq = io_redirect_valid ? 1'h0 : _T_15; // @[IFU.scala 340:21]
  wire [2:0] _T_16 = io_redirect_valid ? 3'h0 : bp1_io_brIdx; // @[IFU.scala 348:29]
  wire [3:0] brIdx = {npcIsSeq,_T_16}; // @[Cat.scala 29:58]
  reg [63:0] _T_19; // @[GTimer.scala 24:20]
  wire [63:0] _T_21 = _T_19 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_23 = pcUpdate & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  wire  _T_25 = ~reset; // @[Debug.scala 56:24]
  wire [42:0] _T_34 = {npcIsSeq,_T_16,npc}; // @[Cat.scala 29:58]
  reg [63:0] _T_39; // @[GTimer.scala 24:20]
  wire [63:0] _T_41 = _T_39 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_43 = _T & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  wire  _T_48 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  reg [63:0] _T_49; // @[GTimer.scala 24:20]
  wire [63:0] _T_51 = _T_49 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_53 = _T_48 & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  wire  _T_62 = ~io_flushVec[0]; // @[IFU.scala 390:41]
  wire  _T_64 = io_imem_resp_ready & io_imem_resp_valid; // @[Decoupled.scala 40:37]
  reg  _T_65; // @[StopWatch.scala 24:20]
  wire  _GEN_3 = io_imem_req_valid | _T_65; // @[StopWatch.scala 30:20]
  wire  _T_66 = |io_flushVec; // @[IFU.scala 393:37]
  BPU_inorder bp1 ( // @[IFU.scala 325:19]
    .clock(bp1_clock),
    .reset(bp1_reset),
    .io_in_pc_valid(bp1_io_in_pc_valid),
    .io_in_pc_bits(bp1_io_in_pc_bits),
    .io_out_target(bp1_io_out_target),
    .io_out_valid(bp1_io_out_valid),
    .io_flush(bp1_io_flush),
    .io_brIdx(bp1_io_brIdx),
    .io_crosslineJump(bp1_io_crosslineJump),
    .MOUFlushICache(bp1_MOUFlushICache),
    .bpuUpdateReq_valid(bp1_bpuUpdateReq_valid),
    .bpuUpdateReq_pc(bp1_bpuUpdateReq_pc),
    .bpuUpdateReq_isMissPredict(bp1_bpuUpdateReq_isMissPredict),
    .bpuUpdateReq_actualTarget(bp1_bpuUpdateReq_actualTarget),
    .bpuUpdateReq_actualTaken(bp1_bpuUpdateReq_actualTaken),
    .bpuUpdateReq_fuOpType(bp1_bpuUpdateReq_fuOpType),
    .bpuUpdateReq_btbType(bp1_bpuUpdateReq_btbType),
    .bpuUpdateReq_isRVC(bp1_bpuUpdateReq_isRVC),
    .DISPLAY_ENABLE(bp1_DISPLAY_ENABLE),
    .MOUFlushTLB(bp1_MOUFlushTLB)
  );
  assign io_imem_req_valid = io_out_ready; // @[IFU.scala 371:21]
  assign io_imem_req_bits_addr = {pc[38:1],1'h0}; // @[SimpleBus.scala 64:15]
  assign io_imem_req_bits_user = {_T_34,pc}; // @[SimpleBus.scala 69:21]
  assign io_imem_resp_ready = io_out_ready | io_flushVec[0]; // @[IFU.scala 373:22]
  assign io_out_valid = io_imem_resp_valid & _T_62; // @[IFU.scala 390:16]
  assign io_out_bits_instr = io_imem_resp_bits_rdata; // @[IFU.scala 383:21]
  assign io_out_bits_pc = io_imem_resp_bits_user[38:0]; // @[IFU.scala 385:20]
  assign io_out_bits_pnpc = io_imem_resp_bits_user[77:39]; // @[IFU.scala 386:22]
  assign io_out_bits_exceptionVec_12 = io_ipf; // @[IFU.scala 389:44]
  assign io_out_bits_brIdx = io_imem_resp_bits_user[81:78]; // @[IFU.scala 387:23]
  assign io_flushVec = io_redirect_valid ? 4'hf : 4'h0; // @[IFU.scala 366:15]
  assign _T_65_0 = _T_65;
  assign _T_66_0 = _T_66;
  assign bp1_clock = clock;
  assign bp1_reset = reset;
  assign bp1_io_in_pc_valid = io_imem_req_ready & io_imem_req_valid; // @[IFU.scala 351:22]
  assign bp1_io_in_pc_bits = io_redirect_valid ? io_redirect_target : _T_12; // @[IFU.scala 352:21]
  assign bp1_io_flush = io_redirect_valid; // @[IFU.scala 357:16]
  assign bp1_MOUFlushICache = flushICache;
  assign bp1_bpuUpdateReq_valid = _T_243_valid;
  assign bp1_bpuUpdateReq_pc = _T_243_pc;
  assign bp1_bpuUpdateReq_isMissPredict = _T_243_isMissPredict;
  assign bp1_bpuUpdateReq_actualTarget = _T_243_actualTarget;
  assign bp1_bpuUpdateReq_actualTaken = _T_243_actualTaken;
  assign bp1_bpuUpdateReq_fuOpType = _T_243_fuOpType;
  assign bp1_bpuUpdateReq_btbType = _T_243_btbType;
  assign bp1_bpuUpdateReq_isRVC = _T_243_isRVC;
  assign bp1_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign bp1_MOUFlushTLB = flushTLB;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  pc = _RAND_0[38:0];
  _RAND_1 = {1{`RANDOM}};
  crosslineJumpLatch = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  crosslineJumpTarget = _RAND_2[38:0];
  _RAND_3 = {2{`RANDOM}};
  _T_19 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  _T_39 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  _T_49 = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  _T_65 = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      pc <= 39'h80000000;
    end else if (pcUpdate) begin
      if (io_redirect_valid) begin
        pc <= io_redirect_target;
      end else if (crosslineJumpLatch) begin
        pc <= crosslineJumpTarget;
      end else if (bp1_io_out_valid) begin
        if (bp1_io_crosslineJump) begin
          if (pc[1]) begin
            pc <= _T_3;
          end else begin
            pc <= _T_5;
          end
        end else begin
          pc <= bp1_io_out_target;
        end
      end else if (pc[1]) begin
        pc <= _T_3;
      end else begin
        pc <= _T_5;
      end
    end
    if (reset) begin
      crosslineJumpLatch <= 1'h0;
    end else if (_T_6) begin
      if (bp1_io_flush) begin
        crosslineJumpLatch <= 1'h0;
      end else begin
        crosslineJumpLatch <= _T_8;
      end
    end
    if (bp1_io_crosslineJump) begin
      crosslineJumpTarget <= bp1_io_out_target;
    end
    if (reset) begin
      _T_19 <= 64'h0;
    end else begin
      _T_19 <= _T_21;
    end
    if (reset) begin
      _T_39 <= 64'h0;
    end else begin
      _T_39 <= _T_41;
    end
    if (reset) begin
      _T_49 <= 64'h0;
    end else begin
      _T_49 <= _T_51;
    end
    if (reset) begin
      _T_65 <= 1'h0;
    end else if (_T_64) begin
      _T_65 <= 1'h0;
    end else begin
      _T_65 <= _GEN_3;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_23 & _T_25) begin
          $fwrite(32'h80000002,"[%d] IFU_inorder: ",_T_19); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_23 & _T_25) begin
          $fwrite(32'h80000002,"[IFUPC] pc:%x pcUpdate:%d npc:%x RedValid:%d RedTarget:%x LJL:%d LJTarget:%x LJ:%d snpc:%x bpValid:%d pnpn:%x \n",pc,pcUpdate,npc,io_redirect_valid,io_redirect_target,crosslineJumpLatch,crosslineJumpTarget,bp1_io_crosslineJump,snpc,bp1_io_out_valid,pnpc); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_43 & _T_25) begin
          $fwrite(32'h80000002,"[%d] IFU_inorder: ",_T_39); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_43 & _T_25) begin
          $fwrite(32'h80000002,"[IFI] pc=%x user=%x %x %x %x \n",io_imem_req_bits_addr,io_imem_req_bits_user,io_redirect_valid,bp1_io_brIdx,brIdx); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_25) begin
          $fwrite(32'h80000002,"[%d] IFU_inorder: ",_T_49); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_53 & _T_25) begin
          $fwrite(32'h80000002,"[IFO] pc=%x inst=%x\n",io_out_bits_pc,io_out_bits_instr); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module NaiveRVCAlignBuffer(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [63:0] io_in_bits_instr,
  input  [38:0] io_in_bits_pc,
  input  [38:0] io_in_bits_pnpc,
  input         io_in_bits_exceptionVec_12,
  input  [3:0]  io_in_bits_brIdx,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_instr,
  output [38:0] io_out_bits_pc,
  output [38:0] io_out_bits_pnpc,
  output        io_out_bits_exceptionVec_12,
  output [3:0]  io_out_bits_brIdx,
  output        io_out_bits_crossPageIPFFix,
  input         io_flush,
  input         DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[NaiveIBF.scala 39:22]
  wire  _T_83 = state == 2'h2; // @[NaiveIBF.scala 90:23]
  wire  _T_84 = state == 2'h3; // @[NaiveIBF.scala 90:47]
  wire  _T_85 = _T_83 | _T_84; // @[NaiveIBF.scala 90:38]
  wire [79:0] instIn = {16'h0,io_in_bits_instr}; // @[Cat.scala 29:58]
  reg [15:0] specialInstR; // @[NaiveIBF.scala 66:25]
  wire [31:0] _T_87 = {instIn[15:0],specialInstR}; // @[Cat.scala 29:58]
  wire  _T_1 = state == 2'h0; // @[NaiveIBF.scala 41:28]
  reg [2:0] pcOffsetR; // @[NaiveIBF.scala 40:26]
  wire [2:0] pcOffset = _T_1 ? io_in_bits_pc[2:0] : pcOffsetR; // @[NaiveIBF.scala 41:21]
  wire  _T_92 = 3'h0 == pcOffset; // @[LookupTree.scala 24:34]
  wire [31:0] _T_96 = _T_92 ? instIn[31:0] : 32'h0; // @[Mux.scala 27:72]
  wire  _T_93 = 3'h2 == pcOffset; // @[LookupTree.scala 24:34]
  wire [31:0] _T_97 = _T_93 ? instIn[47:16] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_100 = _T_96 | _T_97; // @[Mux.scala 27:72]
  wire  _T_94 = 3'h4 == pcOffset; // @[LookupTree.scala 24:34]
  wire [31:0] _T_98 = _T_94 ? instIn[63:32] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_101 = _T_100 | _T_98; // @[Mux.scala 27:72]
  wire  _T_95 = 3'h6 == pcOffset; // @[LookupTree.scala 24:34]
  wire [31:0] _T_99 = _T_95 ? instIn[79:48] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_102 = _T_101 | _T_99; // @[Mux.scala 27:72]
  wire [31:0] instr = _T_85 ? _T_87 : _T_102; // @[NaiveIBF.scala 90:15]
  wire  isRVC = instr[1:0] != 2'h3; // @[NaiveIBF.scala 34:26]
  wire  _T_3 = pcOffset == 3'h0; // @[NaiveIBF.scala 48:28]
  wire  _T_4 = ~isRVC; // @[NaiveIBF.scala 48:40]
  wire  _T_6 = _T_4 | io_in_bits_brIdx[0]; // @[NaiveIBF.scala 48:47]
  wire  _T_7 = _T_3 & _T_6; // @[NaiveIBF.scala 48:36]
  wire  _T_8 = pcOffset == 3'h4; // @[NaiveIBF.scala 48:72]
  wire  _T_12 = _T_8 & _T_6; // @[NaiveIBF.scala 48:80]
  wire  _T_13 = _T_7 | _T_12; // @[NaiveIBF.scala 48:60]
  wire  _T_14 = pcOffset == 3'h2; // @[NaiveIBF.scala 48:116]
  wire  _T_16 = isRVC | io_in_bits_brIdx[1]; // @[NaiveIBF.scala 48:134]
  wire  _T_17 = _T_14 & _T_16; // @[NaiveIBF.scala 48:124]
  wire  _T_18 = _T_13 | _T_17; // @[NaiveIBF.scala 48:104]
  wire  _T_19 = pcOffset == 3'h6; // @[NaiveIBF.scala 48:159]
  wire  _T_20 = _T_19 & isRVC; // @[NaiveIBF.scala 48:167]
  wire  rvcFinish = _T_18 | _T_20; // @[NaiveIBF.scala 48:147]
  wire  _T_23 = ~io_in_bits_brIdx[0]; // @[NaiveIBF.scala 51:47]
  wire  _T_24 = isRVC & _T_23; // @[NaiveIBF.scala 51:44]
  wire  _T_25 = _T_3 & _T_24; // @[NaiveIBF.scala 51:34]
  wire  _T_30 = _T_8 & _T_24; // @[NaiveIBF.scala 51:78]
  wire  _T_31 = _T_25 | _T_30; // @[NaiveIBF.scala 51:58]
  wire  _T_34 = _T_14 & _T_4; // @[NaiveIBF.scala 51:122]
  wire  _T_36 = ~io_in_bits_brIdx[1]; // @[NaiveIBF.scala 51:135]
  wire  _T_37 = _T_34 & _T_36; // @[NaiveIBF.scala 51:132]
  wire  rvcNext = _T_31 | _T_37; // @[NaiveIBF.scala 51:102]
  wire  _T_40 = _T_19 & _T_4; // @[NaiveIBF.scala 52:37]
  wire  _T_42 = ~io_in_bits_brIdx[2]; // @[NaiveIBF.scala 52:50]
  wire  rvcSpecial = _T_40 & _T_42; // @[NaiveIBF.scala 52:47]
  wire  rvcSpecialJump = _T_40 & io_in_bits_brIdx[2]; // @[NaiveIBF.scala 53:51]
  wire  pnpcIsSeq = io_in_bits_brIdx[3]; // @[NaiveIBF.scala 54:24]
  wire  _T_48 = state == 2'h1; // @[NaiveIBF.scala 57:45]
  wire  _T_49 = _T_1 | _T_48; // @[NaiveIBF.scala 57:36]
  wire  _T_50 = _T_49 & rvcSpecial; // @[NaiveIBF.scala 57:58]
  wire  _T_51 = _T_50 & io_in_valid; // @[NaiveIBF.scala 57:72]
  wire  _T_52 = ~pnpcIsSeq; // @[NaiveIBF.scala 57:90]
  wire  flushIFU = _T_51 & _T_52; // @[NaiveIBF.scala 57:87]
  reg [63:0] _T_53; // @[GTimer.scala 24:20]
  wire [63:0] _T_55 = _T_53 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_57 = flushIFU & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  wire  _T_59 = ~reset; // @[Debug.scala 56:24]
  wire  _T_62 = ~flushIFU; // @[NaiveIBF.scala 59:10]
  wire  _T_64 = _T_62 | reset; // @[NaiveIBF.scala 59:9]
  wire  _T_65 = ~_T_64; // @[NaiveIBF.scala 59:9]
  wire  _T_69 = rvcSpecial | rvcSpecialJump; // @[NaiveIBF.scala 60:81]
  wire  _T_70 = _T_49 & _T_69; // @[NaiveIBF.scala 60:66]
  wire  _T_71 = _T_70 & io_in_valid; // @[NaiveIBF.scala 60:100]
  wire  loadNextInstline = _T_71 & pnpcIsSeq; // @[NaiveIBF.scala 60:115]
  reg [38:0] specialPCR; // @[NaiveIBF.scala 64:23]
  reg [38:0] specialNPCR; // @[NaiveIBF.scala 65:24]
  reg  specialIPFR; // @[NaiveIBF.scala 67:28]
  wire  _T_79 = io_in_bits_pnpc[2:0] == 3'h4; // @[NaiveIBF.scala 69:78]
  wire  _T_80 = _T_34 & _T_79; // @[NaiveIBF.scala 69:54]
  wire  rvcForceLoadNext = _T_80 & _T_36; // @[NaiveIBF.scala 69:86]
  wire  _T_105 = ~io_flush; // @[NaiveIBF.scala 97:8]
  wire  _T_106 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_107 = rvcFinish | rvcNext; // @[NaiveIBF.scala 100:28]
  wire  _T_108 = rvcFinish | rvcForceLoadNext; // @[NaiveIBF.scala 101:28]
  wire [38:0] _T_110 = io_in_bits_pc + 39'h2; // @[NaiveIBF.scala 103:76]
  wire [38:0] _T_112 = io_in_bits_pc + 39'h4; // @[NaiveIBF.scala 103:95]
  wire [38:0] _T_113 = isRVC ? _T_110 : _T_112; // @[NaiveIBF.scala 103:55]
  wire [38:0] _T_114 = rvcFinish ? io_in_bits_pnpc : _T_113; // @[NaiveIBF.scala 103:23]
  wire  _T_115 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_116 = _T_115 & rvcFinish; // @[NaiveIBF.scala 104:28]
  wire  _T_118 = _T_115 & rvcNext; // @[NaiveIBF.scala 105:28]
  wire [2:0] _T_119 = isRVC ? 3'h2 : 3'h4; // @[NaiveIBF.scala 107:38]
  wire [2:0] _T_121 = pcOffset + _T_119; // @[NaiveIBF.scala 107:33]
  wire  _T_122 = rvcSpecial & io_in_valid; // @[NaiveIBF.scala 109:25]
  wire  _T_126 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire [38:0] _T_131 = {io_in_bits_pc[38:3],pcOffsetR}; // @[Cat.scala 29:58]
  wire  _T_149 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_153 = 2'h3 == state; // @[Conditional.scala 37:30]
  wire [38:0] _GEN_27 = _T_153 ? specialPCR : 39'h0; // @[Conditional.scala 39:67]
  wire [38:0] _GEN_32 = _T_149 ? specialPCR : _GEN_27; // @[Conditional.scala 39:67]
  wire [38:0] _GEN_40 = _T_126 ? _T_131 : _GEN_32; // @[Conditional.scala 39:67]
  wire [38:0] pcOut = _T_106 ? io_in_bits_pc : _GEN_40; // @[Conditional.scala 40:58]
  wire  _T_124 = rvcSpecialJump & io_in_valid; // @[NaiveIBF.scala 115:29]
  wire [38:0] _T_133 = pcOut + 39'h2; // @[NaiveIBF.scala 127:68]
  wire [38:0] _T_135 = pcOut + 39'h4; // @[NaiveIBF.scala 127:79]
  wire [38:0] _T_136 = isRVC ? _T_133 : _T_135; // @[NaiveIBF.scala 127:55]
  wire [38:0] _T_137 = rvcFinish ? io_in_bits_pnpc : _T_136; // @[NaiveIBF.scala 127:23]
  wire [38:0] _T_151 = specialPCR + 39'h4; // @[NaiveIBF.scala 150:31]
  wire [38:0] _GEN_28 = _T_153 ? specialNPCR : 39'h0; // @[Conditional.scala 39:67]
  wire  _GEN_29 = _T_153 & io_in_valid; // @[Conditional.scala 39:67]
  wire [38:0] _GEN_33 = _T_149 ? _T_151 : _GEN_28; // @[Conditional.scala 39:67]
  wire  _GEN_34 = _T_149 ? io_in_valid : _GEN_29; // @[Conditional.scala 39:67]
  wire  _GEN_35 = _T_149 ? 1'h0 : _T_153; // @[Conditional.scala 39:67]
  wire  _GEN_38 = _T_126 ? _T_107 : _GEN_34; // @[Conditional.scala 39:67]
  wire  _GEN_39 = _T_126 ? _T_108 : _GEN_35; // @[Conditional.scala 39:67]
  wire [38:0] _GEN_41 = _T_126 ? _T_137 : _GEN_33; // @[Conditional.scala 39:67]
  wire  canGo = _T_106 ? _T_107 : _GEN_38; // @[Conditional.scala 40:58]
  wire  canIn = _T_106 ? _T_108 : _GEN_39; // @[Conditional.scala 40:58]
  wire [38:0] pnpcOut = _T_106 ? _T_114 : _GEN_41; // @[Conditional.scala 40:58]
  wire  _T_157 = pnpcOut == _T_135; // @[NaiveIBF.scala 185:37]
  wire  _T_159 = _T_157 & _T_4; // @[NaiveIBF.scala 185:51]
  wire  _T_162 = pnpcOut == _T_133; // @[NaiveIBF.scala 185:74]
  wire  _T_163 = _T_162 & isRVC; // @[NaiveIBF.scala 185:88]
  wire  _T_164 = _T_159 | _T_163; // @[NaiveIBF.scala 185:62]
  wire  _T_165 = _T_164 ? 1'h0 : 1'h1; // @[NaiveIBF.scala 185:27]
  wire  _T_167 = ~io_in_valid; // @[NaiveIBF.scala 188:19]
  wire  _T_169 = _T_115 & canIn; // @[NaiveIBF.scala 188:50]
  wire  _T_170 = _T_167 | _T_169; // @[NaiveIBF.scala 188:32]
  wire  _T_174 = _T_84 | _T_83; // @[NaiveIBF.scala 191:133]
  wire  _T_175 = specialIPFR & _T_174; // @[NaiveIBF.scala 191:102]
  wire  _T_180 = io_in_bits_exceptionVec_12 & _T_174; // @[NaiveIBF.scala 192:74]
  wire  _T_181 = ~specialIPFR; // @[NaiveIBF.scala 192:133]
  assign io_in_ready = _T_170 | loadNextInstline; // @[NaiveIBF.scala 188:15]
  assign io_out_valid = io_in_valid & canGo; // @[NaiveIBF.scala 187:16]
  assign io_out_bits_instr = {{32'd0}, instr}; // @[NaiveIBF.scala 184:21]
  assign io_out_bits_pc = _T_106 ? io_in_bits_pc : _GEN_40; // @[NaiveIBF.scala 182:18]
  assign io_out_bits_pnpc = _T_106 ? _T_114 : _GEN_41; // @[NaiveIBF.scala 183:20]
  assign io_out_bits_exceptionVec_12 = io_in_bits_exceptionVec_12 | _T_175; // @[NaiveIBF.scala 190:28 NaiveIBF.scala 191:44]
  assign io_out_bits_brIdx = {{3'd0}, _T_165}; // @[NaiveIBF.scala 185:21]
  assign io_out_bits_crossPageIPFFix = _T_180 & _T_181; // @[NaiveIBF.scala 192:31]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  specialInstR = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  pcOffsetR = _RAND_2[2:0];
  _RAND_3 = {2{`RANDOM}};
  _T_53 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  specialPCR = _RAND_4[38:0];
  _RAND_5 = {2{`RANDOM}};
  specialNPCR = _RAND_5[38:0];
  _RAND_6 = {1{`RANDOM}};
  specialIPFR = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else if (_T_105) begin
      if (_T_106) begin
        if (_T_124) begin
          state <= 2'h3;
        end else if (_T_122) begin
          state <= 2'h2;
        end else if (_T_118) begin
          state <= 2'h1;
        end else if (_T_116) begin
          state <= 2'h0;
        end
      end else if (_T_126) begin
        if (_T_124) begin
          state <= 2'h3;
        end else if (_T_122) begin
          state <= 2'h2;
        end else if (_T_118) begin
          state <= 2'h1;
        end else if (_T_116) begin
          state <= 2'h0;
        end
      end else if (_T_149) begin
        if (_T_115) begin
          state <= 2'h1;
        end
      end else if (_T_153) begin
        if (_T_115) begin
          state <= 2'h0;
        end
      end
    end else begin
      state <= 2'h0;
    end
    if (_T_105) begin
      if (_T_106) begin
        if (_T_124) begin
          specialInstR <= io_in_bits_instr[63:48];
        end else if (_T_122) begin
          specialInstR <= io_in_bits_instr[63:48];
        end
      end else if (_T_126) begin
        if (_T_124) begin
          specialInstR <= io_in_bits_instr[63:48];
        end else if (_T_122) begin
          specialInstR <= io_in_bits_instr[63:48];
        end
      end
    end
    if (reset) begin
      pcOffsetR <= 3'h0;
    end else if (_T_105) begin
      if (_T_106) begin
        if (_T_118) begin
          pcOffsetR <= _T_121;
        end
      end else if (_T_126) begin
        if (_T_118) begin
          pcOffsetR <= _T_121;
        end
      end else if (_T_149) begin
        if (_T_115) begin
          pcOffsetR <= 3'h2;
        end
      end
    end
    if (reset) begin
      _T_53 <= 64'h0;
    end else begin
      _T_53 <= _T_55;
    end
    if (_T_105) begin
      if (_T_106) begin
        if (_T_124) begin
          if (_T_106) begin
            specialPCR <= io_in_bits_pc;
          end else if (_T_126) begin
            specialPCR <= _T_131;
          end else if (!(_T_149)) begin
            if (!(_T_153)) begin
              specialPCR <= 39'h0;
            end
          end
        end else if (_T_122) begin
          if (_T_106) begin
            specialPCR <= io_in_bits_pc;
          end else if (_T_126) begin
            specialPCR <= _T_131;
          end else if (!(_T_149)) begin
            if (!(_T_153)) begin
              specialPCR <= 39'h0;
            end
          end
        end
      end else if (_T_126) begin
        if (_T_124) begin
          if (_T_106) begin
            specialPCR <= io_in_bits_pc;
          end else if (_T_126) begin
            specialPCR <= _T_131;
          end else if (!(_T_149)) begin
            if (!(_T_153)) begin
              specialPCR <= 39'h0;
            end
          end
        end else if (_T_122) begin
          if (_T_106) begin
            specialPCR <= io_in_bits_pc;
          end else if (_T_126) begin
            specialPCR <= _T_131;
          end else if (!(_T_149)) begin
            if (!(_T_153)) begin
              specialPCR <= 39'h0;
            end
          end
        end
      end
    end
    if (_T_105) begin
      if (_T_106) begin
        if (_T_124) begin
          specialNPCR <= io_in_bits_pnpc;
        end
      end else if (_T_126) begin
        if (_T_124) begin
          specialNPCR <= io_in_bits_pnpc;
        end
      end
    end
    if (reset) begin
      specialIPFR <= 1'h0;
    end else if (_T_105) begin
      if (_T_106) begin
        if (_T_124) begin
          specialIPFR <= io_in_bits_exceptionVec_12;
        end else if (_T_122) begin
          specialIPFR <= io_in_bits_exceptionVec_12;
        end
      end else if (_T_126) begin
        if (_T_124) begin
          specialIPFR <= io_in_bits_exceptionVec_12;
        end else if (_T_122) begin
          specialIPFR <= io_in_bits_exceptionVec_12;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_57 & _T_59) begin
          $fwrite(32'h80000002,"[%d] NaiveRVCAlignBuffer: ",_T_53); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_57 & _T_59) begin
          $fwrite(32'h80000002,"flushIFU at pc %x offset %x\n",io_in_bits_pc,pcOffset); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_65) begin
          $fwrite(32'h80000002,"Assertion failed\n    at NaiveIBF.scala:59 assert(!flushIFU)\n"); // @[NaiveIBF.scala 59:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_65) begin
          $fatal; // @[NaiveIBF.scala 59:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Decoder(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [63:0] io_in_bits_instr,
  input  [38:0] io_in_bits_pc,
  input  [38:0] io_in_bits_pnpc,
  input         io_in_bits_exceptionVec_12,
  input  [3:0]  io_in_bits_brIdx,
  input         io_in_bits_crossPageIPFFix,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_cf_instr,
  output [38:0] io_out_bits_cf_pc,
  output [38:0] io_out_bits_cf_pnpc,
  output        io_out_bits_cf_exceptionVec_1,
  output        io_out_bits_cf_exceptionVec_2,
  output        io_out_bits_cf_exceptionVec_12,
  output        io_out_bits_cf_intrVec_0,
  output        io_out_bits_cf_intrVec_1,
  output        io_out_bits_cf_intrVec_2,
  output        io_out_bits_cf_intrVec_3,
  output        io_out_bits_cf_intrVec_4,
  output        io_out_bits_cf_intrVec_5,
  output        io_out_bits_cf_intrVec_6,
  output        io_out_bits_cf_intrVec_7,
  output        io_out_bits_cf_intrVec_8,
  output        io_out_bits_cf_intrVec_9,
  output        io_out_bits_cf_intrVec_10,
  output        io_out_bits_cf_intrVec_11,
  output [3:0]  io_out_bits_cf_brIdx,
  output        io_out_bits_cf_crossPageIPFFix,
  output [1:0]  io_out_bits_ctrl_src1Type,
  output [1:0]  io_out_bits_ctrl_src2Type,
  output [2:0]  io_out_bits_ctrl_fuType,
  output [6:0]  io_out_bits_ctrl_fuOpType,
  output [4:0]  io_out_bits_ctrl_rfSrc1,
  output [4:0]  io_out_bits_ctrl_rfSrc2,
  output        io_out_bits_ctrl_rfWen,
  output [4:0]  io_out_bits_ctrl_rfDest,
  output        io_out_bits_ctrl_isNutCoreTrap,
  output [63:0] io_out_bits_data_imm,
  output        io_isWFI,
  input         DISPLAY_ENABLE,
  input         DTLBENABLE,
  input  [11:0] intrVecIDU
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] _T = io_in_bits_instr & 64'h707f; // @[Lookup.scala 31:38]
  wire  _T_1 = 64'h13 == _T; // @[Lookup.scala 31:38]
  wire [63:0] _T_2 = io_in_bits_instr & 64'hfc00707f; // @[Lookup.scala 31:38]
  wire  _T_3 = 64'h1013 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_5 = 64'h2013 == _T; // @[Lookup.scala 31:38]
  wire  _T_7 = 64'h3013 == _T; // @[Lookup.scala 31:38]
  wire  _T_9 = 64'h4013 == _T; // @[Lookup.scala 31:38]
  wire  _T_11 = 64'h5013 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_13 = 64'h6013 == _T; // @[Lookup.scala 31:38]
  wire  _T_15 = 64'h7013 == _T; // @[Lookup.scala 31:38]
  wire  _T_17 = 64'h40005013 == _T_2; // @[Lookup.scala 31:38]
  wire [63:0] _T_18 = io_in_bits_instr & 64'hfe00707f; // @[Lookup.scala 31:38]
  wire  _T_19 = 64'h33 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_21 = 64'h1033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_23 = 64'h2033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_25 = 64'h3033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_27 = 64'h4033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_29 = 64'h5033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_31 = 64'h6033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_33 = 64'h7033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_35 = 64'h40000033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_37 = 64'h40005033 == _T_18; // @[Lookup.scala 31:38]
  wire [63:0] _T_38 = io_in_bits_instr & 64'h7f; // @[Lookup.scala 31:38]
  wire  _T_39 = 64'h17 == _T_38; // @[Lookup.scala 31:38]
  wire  _T_41 = 64'h37 == _T_38; // @[Lookup.scala 31:38]
  wire  _T_43 = 64'h6f == _T_38; // @[Lookup.scala 31:38]
  wire  _T_45 = 64'h67 == _T; // @[Lookup.scala 31:38]
  wire  _T_47 = 64'h63 == _T; // @[Lookup.scala 31:38]
  wire  _T_49 = 64'h1063 == _T; // @[Lookup.scala 31:38]
  wire  _T_51 = 64'h4063 == _T; // @[Lookup.scala 31:38]
  wire  _T_53 = 64'h5063 == _T; // @[Lookup.scala 31:38]
  wire  _T_55 = 64'h6063 == _T; // @[Lookup.scala 31:38]
  wire  _T_57 = 64'h7063 == _T; // @[Lookup.scala 31:38]
  wire  _T_59 = 64'h3 == _T; // @[Lookup.scala 31:38]
  wire  _T_61 = 64'h1003 == _T; // @[Lookup.scala 31:38]
  wire  _T_63 = 64'h2003 == _T; // @[Lookup.scala 31:38]
  wire  _T_65 = 64'h4003 == _T; // @[Lookup.scala 31:38]
  wire  _T_67 = 64'h5003 == _T; // @[Lookup.scala 31:38]
  wire  _T_69 = 64'h23 == _T; // @[Lookup.scala 31:38]
  wire  _T_71 = 64'h1023 == _T; // @[Lookup.scala 31:38]
  wire  _T_73 = 64'h2023 == _T; // @[Lookup.scala 31:38]
  wire  _T_75 = 64'h1b == _T; // @[Lookup.scala 31:38]
  wire  _T_77 = 64'h101b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_79 = 64'h501b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_81 = 64'h4000501b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_83 = 64'h103b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_85 = 64'h503b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_87 = 64'h4000503b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_89 = 64'h3b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_91 = 64'h4000003b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_93 = 64'h6003 == _T; // @[Lookup.scala 31:38]
  wire  _T_95 = 64'h3003 == _T; // @[Lookup.scala 31:38]
  wire  _T_97 = 64'h3023 == _T; // @[Lookup.scala 31:38]
  wire  _T_99 = 64'h6b == _T; // @[Lookup.scala 31:38]
  wire  _T_101 = 64'h2000033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_103 = 64'h2001033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_105 = 64'h2002033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_107 = 64'h2003033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_109 = 64'h2004033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_111 = 64'h2005033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_113 = 64'h2006033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_115 = 64'h2007033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_117 = 64'h200003b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_119 = 64'h200403b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_121 = 64'h200503b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_123 = 64'h200603b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_125 = 64'h200703b == _T_18; // @[Lookup.scala 31:38]
  wire [63:0] _T_126 = io_in_bits_instr & 64'hffffffff; // @[Lookup.scala 31:38]
  wire  _T_127 = 64'h0 == _T_126; // @[Lookup.scala 31:38]
  wire [63:0] _T_128 = io_in_bits_instr & 64'he003; // @[Lookup.scala 31:38]
  wire  _T_129 = 64'h0 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_131 = 64'h4000 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_133 = 64'h6000 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_135 = 64'hc000 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_137 = 64'he000 == _T_128; // @[Lookup.scala 31:38]
  wire [63:0] _T_138 = io_in_bits_instr & 64'hef83; // @[Lookup.scala 31:38]
  wire  _T_139 = 64'h1 == _T_138; // @[Lookup.scala 31:38]
  wire  _T_141 = 64'h1 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_143 = 64'h2001 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_145 = 64'h4001 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_147 = 64'h6101 == _T_138; // @[Lookup.scala 31:38]
  wire  _T_149 = 64'h6001 == _T_128; // @[Lookup.scala 31:38]
  wire [63:0] _T_150 = io_in_bits_instr & 64'hec03; // @[Lookup.scala 31:38]
  wire  _T_151 = 64'h8001 == _T_150; // @[Lookup.scala 31:38]
  wire  _T_153 = 64'h8401 == _T_150; // @[Lookup.scala 31:38]
  wire  _T_155 = 64'h8801 == _T_150; // @[Lookup.scala 31:38]
  wire [63:0] _T_156 = io_in_bits_instr & 64'hfc63; // @[Lookup.scala 31:38]
  wire  _T_157 = 64'h8c01 == _T_156; // @[Lookup.scala 31:38]
  wire  _T_159 = 64'h8c21 == _T_156; // @[Lookup.scala 31:38]
  wire  _T_161 = 64'h8c41 == _T_156; // @[Lookup.scala 31:38]
  wire  _T_163 = 64'h8c61 == _T_156; // @[Lookup.scala 31:38]
  wire  _T_165 = 64'h9c01 == _T_156; // @[Lookup.scala 31:38]
  wire  _T_167 = 64'h9c21 == _T_156; // @[Lookup.scala 31:38]
  wire  _T_169 = 64'ha001 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_171 = 64'hc001 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_173 = 64'he001 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_175 = 64'h2 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_177 = 64'h4002 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_179 = 64'h6002 == _T_128; // @[Lookup.scala 31:38]
  wire [63:0] _T_180 = io_in_bits_instr & 64'hf07f; // @[Lookup.scala 31:38]
  wire  _T_181 = 64'h8002 == _T_180; // @[Lookup.scala 31:38]
  wire [63:0] _T_182 = io_in_bits_instr & 64'hf003; // @[Lookup.scala 31:38]
  wire  _T_183 = 64'h8002 == _T_182; // @[Lookup.scala 31:38]
  wire [63:0] _T_184 = io_in_bits_instr & 64'hffff; // @[Lookup.scala 31:38]
  wire  _T_185 = 64'h9002 == _T_184; // @[Lookup.scala 31:38]
  wire  _T_187 = 64'h9002 == _T_180; // @[Lookup.scala 31:38]
  wire  _T_189 = 64'h9002 == _T_182; // @[Lookup.scala 31:38]
  wire  _T_191 = 64'hc002 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_193 = 64'he002 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_195 = 64'h73 == _T_126; // @[Lookup.scala 31:38]
  wire  _T_197 = 64'h100073 == _T_126; // @[Lookup.scala 31:38]
  wire  _T_199 = 64'h30200073 == _T_126; // @[Lookup.scala 31:38]
  wire  _T_201 = 64'hf == _T; // @[Lookup.scala 31:38]
  wire  _T_203 = 64'h10500073 == _T_126; // @[Lookup.scala 31:38]
  wire  _T_205 = 64'h10200073 == _T_126; // @[Lookup.scala 31:38]
  wire [63:0] _T_206 = io_in_bits_instr & 64'hfe007fff; // @[Lookup.scala 31:38]
  wire  _T_207 = 64'h12000073 == _T_206; // @[Lookup.scala 31:38]
  wire [63:0] _T_208 = io_in_bits_instr & 64'hf9f0707f; // @[Lookup.scala 31:38]
  wire  _T_209 = 64'h1000302f == _T_208; // @[Lookup.scala 31:38]
  wire  _T_211 = 64'h1000202f == _T_208; // @[Lookup.scala 31:38]
  wire [63:0] _T_212 = io_in_bits_instr & 64'hf800707f; // @[Lookup.scala 31:38]
  wire  _T_213 = 64'h1800302f == _T_212; // @[Lookup.scala 31:38]
  wire  _T_215 = 64'h1800202f == _T_212; // @[Lookup.scala 31:38]
  wire [63:0] _T_216 = io_in_bits_instr & 64'hf800607f; // @[Lookup.scala 31:38]
  wire  _T_217 = 64'h800202f == _T_216; // @[Lookup.scala 31:38]
  wire  _T_219 = 64'h202f == _T_216; // @[Lookup.scala 31:38]
  wire  _T_221 = 64'h2000202f == _T_216; // @[Lookup.scala 31:38]
  wire  _T_223 = 64'h6000202f == _T_216; // @[Lookup.scala 31:38]
  wire  _T_225 = 64'h4000202f == _T_216; // @[Lookup.scala 31:38]
  wire  _T_227 = 64'h8000202f == _T_216; // @[Lookup.scala 31:38]
  wire  _T_229 = 64'ha000202f == _T_216; // @[Lookup.scala 31:38]
  wire  _T_231 = 64'hc000202f == _T_216; // @[Lookup.scala 31:38]
  wire  _T_233 = 64'he000202f == _T_216; // @[Lookup.scala 31:38]
  wire  _T_235 = 64'h1073 == _T; // @[Lookup.scala 31:38]
  wire  _T_237 = 64'h2073 == _T; // @[Lookup.scala 31:38]
  wire  _T_239 = 64'h3073 == _T; // @[Lookup.scala 31:38]
  wire  _T_241 = 64'h5073 == _T; // @[Lookup.scala 31:38]
  wire  _T_243 = 64'h6073 == _T; // @[Lookup.scala 31:38]
  wire  _T_245 = 64'h7073 == _T; // @[Lookup.scala 31:38]
  wire  _T_247 = 64'h100f == _T_126; // @[Lookup.scala 31:38]
  wire  _T_249 = 64'hb == _T_18; // @[Lookup.scala 31:38]
  wire  _T_251 = 64'h400b == _T_18; // @[Lookup.scala 31:38]
  wire [63:0] _T_252 = io_in_bits_instr & 64'hfff0707f; // @[Lookup.scala 31:38]
  wire  _T_253 = 64'h100b == _T_252; // @[Lookup.scala 31:38]
  wire  _T_255 = 64'h200100b == _T_252; // @[Lookup.scala 31:38]
  wire  _T_257 = 64'h400100b == _T_252; // @[Lookup.scala 31:38]
  wire  _T_259 = 64'h600100b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_261 = 64'h800100b == _T_252; // @[Lookup.scala 31:38]
  wire  _T_263 = 64'h200b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_265 = 64'h300b == _T; // @[Lookup.scala 31:38]
  wire  _T_267 = 64'h500b == _T; // @[Lookup.scala 31:38]
  wire  _T_269 = 64'h600b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_271 = 64'h700b == _T; // @[Lookup.scala 31:38]
  wire [4:0] _T_272 = _T_271 ? 5'h17 : 5'h0; // @[Lookup.scala 33:37]
  wire [4:0] _T_273 = _T_269 ? 5'h16 : _T_272; // @[Lookup.scala 33:37]
  wire [4:0] _T_274 = _T_267 ? 5'h15 : _T_273; // @[Lookup.scala 33:37]
  wire [4:0] _T_275 = _T_265 ? 5'h10 : _T_274; // @[Lookup.scala 33:37]
  wire [4:0] _T_276 = _T_263 ? 5'h16 : _T_275; // @[Lookup.scala 33:37]
  wire [4:0] _T_277 = _T_261 ? 5'h16 : _T_276; // @[Lookup.scala 33:37]
  wire [4:0] _T_278 = _T_259 ? 5'h16 : _T_277; // @[Lookup.scala 33:37]
  wire [4:0] _T_279 = _T_257 ? 5'h1f : _T_278; // @[Lookup.scala 33:37]
  wire [4:0] _T_280 = _T_255 ? 5'h16 : _T_279; // @[Lookup.scala 33:37]
  wire [4:0] _T_281 = _T_253 ? 5'h16 : _T_280; // @[Lookup.scala 33:37]
  wire [4:0] _T_282 = _T_251 ? 5'h16 : _T_281; // @[Lookup.scala 33:37]
  wire [4:0] _T_283 = _T_249 ? 5'h16 : _T_282; // @[Lookup.scala 33:37]
  wire [4:0] _T_284 = _T_247 ? 5'h1 : _T_283; // @[Lookup.scala 33:37]
  wire [4:0] _T_285 = _T_245 ? 5'h4 : _T_284; // @[Lookup.scala 33:37]
  wire [4:0] _T_286 = _T_243 ? 5'h4 : _T_285; // @[Lookup.scala 33:37]
  wire [4:0] _T_287 = _T_241 ? 5'h4 : _T_286; // @[Lookup.scala 33:37]
  wire [4:0] _T_288 = _T_239 ? 5'h4 : _T_287; // @[Lookup.scala 33:37]
  wire [4:0] _T_289 = _T_237 ? 5'h4 : _T_288; // @[Lookup.scala 33:37]
  wire [4:0] _T_290 = _T_235 ? 5'h4 : _T_289; // @[Lookup.scala 33:37]
  wire [4:0] _T_291 = _T_233 ? 5'h5 : _T_290; // @[Lookup.scala 33:37]
  wire [4:0] _T_292 = _T_231 ? 5'h5 : _T_291; // @[Lookup.scala 33:37]
  wire [4:0] _T_293 = _T_229 ? 5'h5 : _T_292; // @[Lookup.scala 33:37]
  wire [4:0] _T_294 = _T_227 ? 5'h5 : _T_293; // @[Lookup.scala 33:37]
  wire [4:0] _T_295 = _T_225 ? 5'h5 : _T_294; // @[Lookup.scala 33:37]
  wire [4:0] _T_296 = _T_223 ? 5'h5 : _T_295; // @[Lookup.scala 33:37]
  wire [4:0] _T_297 = _T_221 ? 5'h5 : _T_296; // @[Lookup.scala 33:37]
  wire [4:0] _T_298 = _T_219 ? 5'h5 : _T_297; // @[Lookup.scala 33:37]
  wire [4:0] _T_299 = _T_217 ? 5'h5 : _T_298; // @[Lookup.scala 33:37]
  wire [4:0] _T_300 = _T_215 ? 5'hf : _T_299; // @[Lookup.scala 33:37]
  wire [4:0] _T_301 = _T_213 ? 5'hf : _T_300; // @[Lookup.scala 33:37]
  wire [4:0] _T_302 = _T_211 ? 5'h4 : _T_301; // @[Lookup.scala 33:37]
  wire [4:0] _T_303 = _T_209 ? 5'h4 : _T_302; // @[Lookup.scala 33:37]
  wire [4:0] _T_304 = _T_207 ? 5'h5 : _T_303; // @[Lookup.scala 33:37]
  wire [4:0] _T_305 = _T_205 ? 5'h4 : _T_304; // @[Lookup.scala 33:37]
  wire [4:0] _T_306 = _T_203 ? 5'h4 : _T_305; // @[Lookup.scala 33:37]
  wire [4:0] _T_307 = _T_201 ? 5'h2 : _T_306; // @[Lookup.scala 33:37]
  wire [4:0] _T_308 = _T_199 ? 5'h4 : _T_307; // @[Lookup.scala 33:37]
  wire [4:0] _T_309 = _T_197 ? 5'h4 : _T_308; // @[Lookup.scala 33:37]
  wire [4:0] _T_310 = _T_195 ? 5'h4 : _T_309; // @[Lookup.scala 33:37]
  wire [4:0] _T_311 = _T_193 ? 5'h2 : _T_310; // @[Lookup.scala 33:37]
  wire [4:0] _T_312 = _T_191 ? 5'h2 : _T_311; // @[Lookup.scala 33:37]
  wire [4:0] _T_313 = _T_189 ? 5'h5 : _T_312; // @[Lookup.scala 33:37]
  wire [4:0] _T_314 = _T_187 ? 5'h4 : _T_313; // @[Lookup.scala 33:37]
  wire [4:0] _T_315 = _T_185 ? 5'h4 : _T_314; // @[Lookup.scala 33:37]
  wire [4:0] _T_316 = _T_183 ? 5'h5 : _T_315; // @[Lookup.scala 33:37]
  wire [4:0] _T_317 = _T_181 ? 5'h4 : _T_316; // @[Lookup.scala 33:37]
  wire [4:0] _T_318 = _T_179 ? 5'h4 : _T_317; // @[Lookup.scala 33:37]
  wire [4:0] _T_319 = _T_177 ? 5'h4 : _T_318; // @[Lookup.scala 33:37]
  wire [4:0] _T_320 = _T_175 ? 5'h4 : _T_319; // @[Lookup.scala 33:37]
  wire [4:0] _T_321 = _T_173 ? 5'h1 : _T_320; // @[Lookup.scala 33:37]
  wire [4:0] _T_322 = _T_171 ? 5'h1 : _T_321; // @[Lookup.scala 33:37]
  wire [4:0] _T_323 = _T_169 ? 5'h7 : _T_322; // @[Lookup.scala 33:37]
  wire [4:0] _T_324 = _T_167 ? 5'h5 : _T_323; // @[Lookup.scala 33:37]
  wire [4:0] _T_325 = _T_165 ? 5'h5 : _T_324; // @[Lookup.scala 33:37]
  wire [4:0] _T_326 = _T_163 ? 5'h5 : _T_325; // @[Lookup.scala 33:37]
  wire [4:0] _T_327 = _T_161 ? 5'h5 : _T_326; // @[Lookup.scala 33:37]
  wire [4:0] _T_328 = _T_159 ? 5'h5 : _T_327; // @[Lookup.scala 33:37]
  wire [4:0] _T_329 = _T_157 ? 5'h5 : _T_328; // @[Lookup.scala 33:37]
  wire [4:0] _T_330 = _T_155 ? 5'h4 : _T_329; // @[Lookup.scala 33:37]
  wire [4:0] _T_331 = _T_153 ? 5'h4 : _T_330; // @[Lookup.scala 33:37]
  wire [4:0] _T_332 = _T_151 ? 5'h4 : _T_331; // @[Lookup.scala 33:37]
  wire [4:0] _T_333 = _T_149 ? 5'h4 : _T_332; // @[Lookup.scala 33:37]
  wire [4:0] _T_334 = _T_147 ? 5'h4 : _T_333; // @[Lookup.scala 33:37]
  wire [4:0] _T_335 = _T_145 ? 5'h4 : _T_334; // @[Lookup.scala 33:37]
  wire [4:0] _T_336 = _T_143 ? 5'h4 : _T_335; // @[Lookup.scala 33:37]
  wire [4:0] _T_337 = _T_141 ? 5'h4 : _T_336; // @[Lookup.scala 33:37]
  wire [4:0] _T_338 = _T_139 ? 5'h4 : _T_337; // @[Lookup.scala 33:37]
  wire [4:0] _T_339 = _T_137 ? 5'h2 : _T_338; // @[Lookup.scala 33:37]
  wire [4:0] _T_340 = _T_135 ? 5'h2 : _T_339; // @[Lookup.scala 33:37]
  wire [4:0] _T_341 = _T_133 ? 5'h4 : _T_340; // @[Lookup.scala 33:37]
  wire [4:0] _T_342 = _T_131 ? 5'h4 : _T_341; // @[Lookup.scala 33:37]
  wire [4:0] _T_343 = _T_129 ? 5'h4 : _T_342; // @[Lookup.scala 33:37]
  wire [4:0] _T_344 = _T_127 ? 5'h0 : _T_343; // @[Lookup.scala 33:37]
  wire [4:0] _T_345 = _T_125 ? 5'h5 : _T_344; // @[Lookup.scala 33:37]
  wire [4:0] _T_346 = _T_123 ? 5'h5 : _T_345; // @[Lookup.scala 33:37]
  wire [4:0] _T_347 = _T_121 ? 5'h5 : _T_346; // @[Lookup.scala 33:37]
  wire [4:0] _T_348 = _T_119 ? 5'h5 : _T_347; // @[Lookup.scala 33:37]
  wire [4:0] _T_349 = _T_117 ? 5'h5 : _T_348; // @[Lookup.scala 33:37]
  wire [4:0] _T_350 = _T_115 ? 5'h5 : _T_349; // @[Lookup.scala 33:37]
  wire [4:0] _T_351 = _T_113 ? 5'h5 : _T_350; // @[Lookup.scala 33:37]
  wire [4:0] _T_352 = _T_111 ? 5'h5 : _T_351; // @[Lookup.scala 33:37]
  wire [4:0] _T_353 = _T_109 ? 5'h5 : _T_352; // @[Lookup.scala 33:37]
  wire [4:0] _T_354 = _T_107 ? 5'h5 : _T_353; // @[Lookup.scala 33:37]
  wire [4:0] _T_355 = _T_105 ? 5'h5 : _T_354; // @[Lookup.scala 33:37]
  wire [4:0] _T_356 = _T_103 ? 5'h5 : _T_355; // @[Lookup.scala 33:37]
  wire [4:0] _T_357 = _T_101 ? 5'h5 : _T_356; // @[Lookup.scala 33:37]
  wire [4:0] _T_358 = _T_99 ? 5'h4 : _T_357; // @[Lookup.scala 33:37]
  wire [4:0] _T_359 = _T_97 ? 5'h2 : _T_358; // @[Lookup.scala 33:37]
  wire [4:0] _T_360 = _T_95 ? 5'h4 : _T_359; // @[Lookup.scala 33:37]
  wire [4:0] _T_361 = _T_93 ? 5'h4 : _T_360; // @[Lookup.scala 33:37]
  wire [4:0] _T_362 = _T_91 ? 5'h5 : _T_361; // @[Lookup.scala 33:37]
  wire [4:0] _T_363 = _T_89 ? 5'h5 : _T_362; // @[Lookup.scala 33:37]
  wire [4:0] _T_364 = _T_87 ? 5'h5 : _T_363; // @[Lookup.scala 33:37]
  wire [4:0] _T_365 = _T_85 ? 5'h5 : _T_364; // @[Lookup.scala 33:37]
  wire [4:0] _T_366 = _T_83 ? 5'h5 : _T_365; // @[Lookup.scala 33:37]
  wire [4:0] _T_367 = _T_81 ? 5'h4 : _T_366; // @[Lookup.scala 33:37]
  wire [4:0] _T_368 = _T_79 ? 5'h4 : _T_367; // @[Lookup.scala 33:37]
  wire [4:0] _T_369 = _T_77 ? 5'h4 : _T_368; // @[Lookup.scala 33:37]
  wire [4:0] _T_370 = _T_75 ? 5'h4 : _T_369; // @[Lookup.scala 33:37]
  wire [4:0] _T_371 = _T_73 ? 5'h2 : _T_370; // @[Lookup.scala 33:37]
  wire [4:0] _T_372 = _T_71 ? 5'h2 : _T_371; // @[Lookup.scala 33:37]
  wire [4:0] _T_373 = _T_69 ? 5'h2 : _T_372; // @[Lookup.scala 33:37]
  wire [4:0] _T_374 = _T_67 ? 5'h4 : _T_373; // @[Lookup.scala 33:37]
  wire [4:0] _T_375 = _T_65 ? 5'h4 : _T_374; // @[Lookup.scala 33:37]
  wire [4:0] _T_376 = _T_63 ? 5'h4 : _T_375; // @[Lookup.scala 33:37]
  wire [4:0] _T_377 = _T_61 ? 5'h4 : _T_376; // @[Lookup.scala 33:37]
  wire [4:0] _T_378 = _T_59 ? 5'h4 : _T_377; // @[Lookup.scala 33:37]
  wire [4:0] _T_379 = _T_57 ? 5'h1 : _T_378; // @[Lookup.scala 33:37]
  wire [4:0] _T_380 = _T_55 ? 5'h1 : _T_379; // @[Lookup.scala 33:37]
  wire [4:0] _T_381 = _T_53 ? 5'h1 : _T_380; // @[Lookup.scala 33:37]
  wire [4:0] _T_382 = _T_51 ? 5'h1 : _T_381; // @[Lookup.scala 33:37]
  wire [4:0] _T_383 = _T_49 ? 5'h1 : _T_382; // @[Lookup.scala 33:37]
  wire [4:0] _T_384 = _T_47 ? 5'h1 : _T_383; // @[Lookup.scala 33:37]
  wire [4:0] _T_385 = _T_45 ? 5'h4 : _T_384; // @[Lookup.scala 33:37]
  wire [4:0] _T_386 = _T_43 ? 5'h7 : _T_385; // @[Lookup.scala 33:37]
  wire [4:0] _T_387 = _T_41 ? 5'h6 : _T_386; // @[Lookup.scala 33:37]
  wire [4:0] _T_388 = _T_39 ? 5'h6 : _T_387; // @[Lookup.scala 33:37]
  wire [4:0] _T_389 = _T_37 ? 5'h5 : _T_388; // @[Lookup.scala 33:37]
  wire [4:0] _T_390 = _T_35 ? 5'h5 : _T_389; // @[Lookup.scala 33:37]
  wire [4:0] _T_391 = _T_33 ? 5'h5 : _T_390; // @[Lookup.scala 33:37]
  wire [4:0] _T_392 = _T_31 ? 5'h5 : _T_391; // @[Lookup.scala 33:37]
  wire [4:0] _T_393 = _T_29 ? 5'h5 : _T_392; // @[Lookup.scala 33:37]
  wire [4:0] _T_394 = _T_27 ? 5'h5 : _T_393; // @[Lookup.scala 33:37]
  wire [4:0] _T_395 = _T_25 ? 5'h5 : _T_394; // @[Lookup.scala 33:37]
  wire [4:0] _T_396 = _T_23 ? 5'h5 : _T_395; // @[Lookup.scala 33:37]
  wire [4:0] _T_397 = _T_21 ? 5'h5 : _T_396; // @[Lookup.scala 33:37]
  wire [4:0] _T_398 = _T_19 ? 5'h5 : _T_397; // @[Lookup.scala 33:37]
  wire [4:0] _T_399 = _T_17 ? 5'h4 : _T_398; // @[Lookup.scala 33:37]
  wire [4:0] _T_400 = _T_15 ? 5'h4 : _T_399; // @[Lookup.scala 33:37]
  wire [4:0] _T_401 = _T_13 ? 5'h4 : _T_400; // @[Lookup.scala 33:37]
  wire [4:0] _T_402 = _T_11 ? 5'h4 : _T_401; // @[Lookup.scala 33:37]
  wire [4:0] _T_403 = _T_9 ? 5'h4 : _T_402; // @[Lookup.scala 33:37]
  wire [4:0] _T_404 = _T_7 ? 5'h4 : _T_403; // @[Lookup.scala 33:37]
  wire [4:0] _T_405 = _T_5 ? 5'h4 : _T_404; // @[Lookup.scala 33:37]
  wire [4:0] _T_406 = _T_3 ? 5'h4 : _T_405; // @[Lookup.scala 33:37]
  wire [4:0] decodeList_0 = _T_1 ? 5'h4 : _T_406; // @[Lookup.scala 33:37]
  wire [2:0] _T_407 = _T_271 ? 3'h5 : 3'h3; // @[Lookup.scala 33:37]
  wire [2:0] _T_408 = _T_269 ? 3'h5 : _T_407; // @[Lookup.scala 33:37]
  wire [2:0] _T_409 = _T_267 ? 3'h1 : _T_408; // @[Lookup.scala 33:37]
  wire [2:0] _T_410 = _T_265 ? 3'h1 : _T_409; // @[Lookup.scala 33:37]
  wire [2:0] _T_411 = _T_263 ? 3'h5 : _T_410; // @[Lookup.scala 33:37]
  wire [2:0] _T_412 = _T_261 ? 3'h5 : _T_411; // @[Lookup.scala 33:37]
  wire [2:0] _T_413 = _T_259 ? 3'h5 : _T_412; // @[Lookup.scala 33:37]
  wire [2:0] _T_414 = _T_257 ? 3'h5 : _T_413; // @[Lookup.scala 33:37]
  wire [2:0] _T_415 = _T_255 ? 3'h5 : _T_414; // @[Lookup.scala 33:37]
  wire [2:0] _T_416 = _T_253 ? 3'h5 : _T_415; // @[Lookup.scala 33:37]
  wire [2:0] _T_417 = _T_251 ? 3'h5 : _T_416; // @[Lookup.scala 33:37]
  wire [2:0] _T_418 = _T_249 ? 3'h5 : _T_417; // @[Lookup.scala 33:37]
  wire [2:0] _T_419 = _T_247 ? 3'h4 : _T_418; // @[Lookup.scala 33:37]
  wire [2:0] _T_420 = _T_245 ? 3'h3 : _T_419; // @[Lookup.scala 33:37]
  wire [2:0] _T_421 = _T_243 ? 3'h3 : _T_420; // @[Lookup.scala 33:37]
  wire [2:0] _T_422 = _T_241 ? 3'h3 : _T_421; // @[Lookup.scala 33:37]
  wire [2:0] _T_423 = _T_239 ? 3'h3 : _T_422; // @[Lookup.scala 33:37]
  wire [2:0] _T_424 = _T_237 ? 3'h3 : _T_423; // @[Lookup.scala 33:37]
  wire [2:0] _T_425 = _T_235 ? 3'h3 : _T_424; // @[Lookup.scala 33:37]
  wire [2:0] _T_426 = _T_233 ? 3'h1 : _T_425; // @[Lookup.scala 33:37]
  wire [2:0] _T_427 = _T_231 ? 3'h1 : _T_426; // @[Lookup.scala 33:37]
  wire [2:0] _T_428 = _T_229 ? 3'h1 : _T_427; // @[Lookup.scala 33:37]
  wire [2:0] _T_429 = _T_227 ? 3'h1 : _T_428; // @[Lookup.scala 33:37]
  wire [2:0] _T_430 = _T_225 ? 3'h1 : _T_429; // @[Lookup.scala 33:37]
  wire [2:0] _T_431 = _T_223 ? 3'h1 : _T_430; // @[Lookup.scala 33:37]
  wire [2:0] _T_432 = _T_221 ? 3'h1 : _T_431; // @[Lookup.scala 33:37]
  wire [2:0] _T_433 = _T_219 ? 3'h1 : _T_432; // @[Lookup.scala 33:37]
  wire [2:0] _T_434 = _T_217 ? 3'h1 : _T_433; // @[Lookup.scala 33:37]
  wire [2:0] _T_435 = _T_215 ? 3'h1 : _T_434; // @[Lookup.scala 33:37]
  wire [2:0] _T_436 = _T_213 ? 3'h1 : _T_435; // @[Lookup.scala 33:37]
  wire [2:0] _T_437 = _T_211 ? 3'h1 : _T_436; // @[Lookup.scala 33:37]
  wire [2:0] _T_438 = _T_209 ? 3'h1 : _T_437; // @[Lookup.scala 33:37]
  wire [2:0] _T_439 = _T_207 ? 3'h4 : _T_438; // @[Lookup.scala 33:37]
  wire [2:0] _T_440 = _T_205 ? 3'h3 : _T_439; // @[Lookup.scala 33:37]
  wire [2:0] _T_441 = _T_203 ? 3'h0 : _T_440; // @[Lookup.scala 33:37]
  wire [2:0] _T_442 = _T_201 ? 3'h4 : _T_441; // @[Lookup.scala 33:37]
  wire [2:0] _T_443 = _T_199 ? 3'h3 : _T_442; // @[Lookup.scala 33:37]
  wire [2:0] _T_444 = _T_197 ? 3'h3 : _T_443; // @[Lookup.scala 33:37]
  wire [2:0] _T_445 = _T_195 ? 3'h3 : _T_444; // @[Lookup.scala 33:37]
  wire [2:0] _T_446 = _T_193 ? 3'h1 : _T_445; // @[Lookup.scala 33:37]
  wire [2:0] _T_447 = _T_191 ? 3'h1 : _T_446; // @[Lookup.scala 33:37]
  wire [2:0] _T_448 = _T_189 ? 3'h0 : _T_447; // @[Lookup.scala 33:37]
  wire [2:0] _T_449 = _T_187 ? 3'h0 : _T_448; // @[Lookup.scala 33:37]
  wire [2:0] _T_450 = _T_185 ? 3'h3 : _T_449; // @[Lookup.scala 33:37]
  wire [2:0] _T_451 = _T_183 ? 3'h0 : _T_450; // @[Lookup.scala 33:37]
  wire [2:0] _T_452 = _T_181 ? 3'h0 : _T_451; // @[Lookup.scala 33:37]
  wire [2:0] _T_453 = _T_179 ? 3'h1 : _T_452; // @[Lookup.scala 33:37]
  wire [2:0] _T_454 = _T_177 ? 3'h1 : _T_453; // @[Lookup.scala 33:37]
  wire [2:0] _T_455 = _T_175 ? 3'h0 : _T_454; // @[Lookup.scala 33:37]
  wire [2:0] _T_456 = _T_173 ? 3'h0 : _T_455; // @[Lookup.scala 33:37]
  wire [2:0] _T_457 = _T_171 ? 3'h0 : _T_456; // @[Lookup.scala 33:37]
  wire [2:0] _T_458 = _T_169 ? 3'h0 : _T_457; // @[Lookup.scala 33:37]
  wire [2:0] _T_459 = _T_167 ? 3'h0 : _T_458; // @[Lookup.scala 33:37]
  wire [2:0] _T_460 = _T_165 ? 3'h0 : _T_459; // @[Lookup.scala 33:37]
  wire [2:0] _T_461 = _T_163 ? 3'h0 : _T_460; // @[Lookup.scala 33:37]
  wire [2:0] _T_462 = _T_161 ? 3'h0 : _T_461; // @[Lookup.scala 33:37]
  wire [2:0] _T_463 = _T_159 ? 3'h0 : _T_462; // @[Lookup.scala 33:37]
  wire [2:0] _T_464 = _T_157 ? 3'h0 : _T_463; // @[Lookup.scala 33:37]
  wire [2:0] _T_465 = _T_155 ? 3'h0 : _T_464; // @[Lookup.scala 33:37]
  wire [2:0] _T_466 = _T_153 ? 3'h0 : _T_465; // @[Lookup.scala 33:37]
  wire [2:0] _T_467 = _T_151 ? 3'h0 : _T_466; // @[Lookup.scala 33:37]
  wire [2:0] _T_468 = _T_149 ? 3'h0 : _T_467; // @[Lookup.scala 33:37]
  wire [2:0] _T_469 = _T_147 ? 3'h0 : _T_468; // @[Lookup.scala 33:37]
  wire [2:0] _T_470 = _T_145 ? 3'h0 : _T_469; // @[Lookup.scala 33:37]
  wire [2:0] _T_471 = _T_143 ? 3'h0 : _T_470; // @[Lookup.scala 33:37]
  wire [2:0] _T_472 = _T_141 ? 3'h0 : _T_471; // @[Lookup.scala 33:37]
  wire [2:0] _T_473 = _T_139 ? 3'h0 : _T_472; // @[Lookup.scala 33:37]
  wire [2:0] _T_474 = _T_137 ? 3'h1 : _T_473; // @[Lookup.scala 33:37]
  wire [2:0] _T_475 = _T_135 ? 3'h1 : _T_474; // @[Lookup.scala 33:37]
  wire [2:0] _T_476 = _T_133 ? 3'h1 : _T_475; // @[Lookup.scala 33:37]
  wire [2:0] _T_477 = _T_131 ? 3'h1 : _T_476; // @[Lookup.scala 33:37]
  wire [2:0] _T_478 = _T_129 ? 3'h0 : _T_477; // @[Lookup.scala 33:37]
  wire [2:0] _T_479 = _T_127 ? 3'h3 : _T_478; // @[Lookup.scala 33:37]
  wire [2:0] _T_480 = _T_125 ? 3'h2 : _T_479; // @[Lookup.scala 33:37]
  wire [2:0] _T_481 = _T_123 ? 3'h2 : _T_480; // @[Lookup.scala 33:37]
  wire [2:0] _T_482 = _T_121 ? 3'h2 : _T_481; // @[Lookup.scala 33:37]
  wire [2:0] _T_483 = _T_119 ? 3'h2 : _T_482; // @[Lookup.scala 33:37]
  wire [2:0] _T_484 = _T_117 ? 3'h2 : _T_483; // @[Lookup.scala 33:37]
  wire [2:0] _T_485 = _T_115 ? 3'h2 : _T_484; // @[Lookup.scala 33:37]
  wire [2:0] _T_486 = _T_113 ? 3'h2 : _T_485; // @[Lookup.scala 33:37]
  wire [2:0] _T_487 = _T_111 ? 3'h2 : _T_486; // @[Lookup.scala 33:37]
  wire [2:0] _T_488 = _T_109 ? 3'h2 : _T_487; // @[Lookup.scala 33:37]
  wire [2:0] _T_489 = _T_107 ? 3'h2 : _T_488; // @[Lookup.scala 33:37]
  wire [2:0] _T_490 = _T_105 ? 3'h2 : _T_489; // @[Lookup.scala 33:37]
  wire [2:0] _T_491 = _T_103 ? 3'h2 : _T_490; // @[Lookup.scala 33:37]
  wire [2:0] _T_492 = _T_101 ? 3'h2 : _T_491; // @[Lookup.scala 33:37]
  wire [2:0] _T_493 = _T_99 ? 3'h3 : _T_492; // @[Lookup.scala 33:37]
  wire [2:0] _T_494 = _T_97 ? 3'h1 : _T_493; // @[Lookup.scala 33:37]
  wire [2:0] _T_495 = _T_95 ? 3'h1 : _T_494; // @[Lookup.scala 33:37]
  wire [2:0] _T_496 = _T_93 ? 3'h1 : _T_495; // @[Lookup.scala 33:37]
  wire [2:0] _T_497 = _T_91 ? 3'h0 : _T_496; // @[Lookup.scala 33:37]
  wire [2:0] _T_498 = _T_89 ? 3'h0 : _T_497; // @[Lookup.scala 33:37]
  wire [2:0] _T_499 = _T_87 ? 3'h0 : _T_498; // @[Lookup.scala 33:37]
  wire [2:0] _T_500 = _T_85 ? 3'h0 : _T_499; // @[Lookup.scala 33:37]
  wire [2:0] _T_501 = _T_83 ? 3'h0 : _T_500; // @[Lookup.scala 33:37]
  wire [2:0] _T_502 = _T_81 ? 3'h0 : _T_501; // @[Lookup.scala 33:37]
  wire [2:0] _T_503 = _T_79 ? 3'h0 : _T_502; // @[Lookup.scala 33:37]
  wire [2:0] _T_504 = _T_77 ? 3'h0 : _T_503; // @[Lookup.scala 33:37]
  wire [2:0] _T_505 = _T_75 ? 3'h0 : _T_504; // @[Lookup.scala 33:37]
  wire [2:0] _T_506 = _T_73 ? 3'h1 : _T_505; // @[Lookup.scala 33:37]
  wire [2:0] _T_507 = _T_71 ? 3'h1 : _T_506; // @[Lookup.scala 33:37]
  wire [2:0] _T_508 = _T_69 ? 3'h1 : _T_507; // @[Lookup.scala 33:37]
  wire [2:0] _T_509 = _T_67 ? 3'h1 : _T_508; // @[Lookup.scala 33:37]
  wire [2:0] _T_510 = _T_65 ? 3'h1 : _T_509; // @[Lookup.scala 33:37]
  wire [2:0] _T_511 = _T_63 ? 3'h1 : _T_510; // @[Lookup.scala 33:37]
  wire [2:0] _T_512 = _T_61 ? 3'h1 : _T_511; // @[Lookup.scala 33:37]
  wire [2:0] _T_513 = _T_59 ? 3'h1 : _T_512; // @[Lookup.scala 33:37]
  wire [2:0] _T_514 = _T_57 ? 3'h0 : _T_513; // @[Lookup.scala 33:37]
  wire [2:0] _T_515 = _T_55 ? 3'h0 : _T_514; // @[Lookup.scala 33:37]
  wire [2:0] _T_516 = _T_53 ? 3'h0 : _T_515; // @[Lookup.scala 33:37]
  wire [2:0] _T_517 = _T_51 ? 3'h0 : _T_516; // @[Lookup.scala 33:37]
  wire [2:0] _T_518 = _T_49 ? 3'h0 : _T_517; // @[Lookup.scala 33:37]
  wire [2:0] _T_519 = _T_47 ? 3'h0 : _T_518; // @[Lookup.scala 33:37]
  wire [2:0] _T_520 = _T_45 ? 3'h0 : _T_519; // @[Lookup.scala 33:37]
  wire [2:0] _T_521 = _T_43 ? 3'h0 : _T_520; // @[Lookup.scala 33:37]
  wire [2:0] _T_522 = _T_41 ? 3'h0 : _T_521; // @[Lookup.scala 33:37]
  wire [2:0] _T_523 = _T_39 ? 3'h0 : _T_522; // @[Lookup.scala 33:37]
  wire [2:0] _T_524 = _T_37 ? 3'h0 : _T_523; // @[Lookup.scala 33:37]
  wire [2:0] _T_525 = _T_35 ? 3'h0 : _T_524; // @[Lookup.scala 33:37]
  wire [2:0] _T_526 = _T_33 ? 3'h0 : _T_525; // @[Lookup.scala 33:37]
  wire [2:0] _T_527 = _T_31 ? 3'h0 : _T_526; // @[Lookup.scala 33:37]
  wire [2:0] _T_528 = _T_29 ? 3'h0 : _T_527; // @[Lookup.scala 33:37]
  wire [2:0] _T_529 = _T_27 ? 3'h0 : _T_528; // @[Lookup.scala 33:37]
  wire [2:0] _T_530 = _T_25 ? 3'h0 : _T_529; // @[Lookup.scala 33:37]
  wire [2:0] _T_531 = _T_23 ? 3'h0 : _T_530; // @[Lookup.scala 33:37]
  wire [2:0] _T_532 = _T_21 ? 3'h0 : _T_531; // @[Lookup.scala 33:37]
  wire [2:0] _T_533 = _T_19 ? 3'h0 : _T_532; // @[Lookup.scala 33:37]
  wire [2:0] _T_534 = _T_17 ? 3'h0 : _T_533; // @[Lookup.scala 33:37]
  wire [2:0] _T_535 = _T_15 ? 3'h0 : _T_534; // @[Lookup.scala 33:37]
  wire [2:0] _T_536 = _T_13 ? 3'h0 : _T_535; // @[Lookup.scala 33:37]
  wire [2:0] _T_537 = _T_11 ? 3'h0 : _T_536; // @[Lookup.scala 33:37]
  wire [2:0] _T_538 = _T_9 ? 3'h0 : _T_537; // @[Lookup.scala 33:37]
  wire [2:0] _T_539 = _T_7 ? 3'h0 : _T_538; // @[Lookup.scala 33:37]
  wire [2:0] _T_540 = _T_5 ? 3'h0 : _T_539; // @[Lookup.scala 33:37]
  wire [2:0] _T_541 = _T_3 ? 3'h0 : _T_540; // @[Lookup.scala 33:37]
  wire [2:0] decodeList_1 = _T_1 ? 3'h0 : _T_541; // @[Lookup.scala 33:37]
  wire [3:0] _T_542 = _T_271 ? 4'he : 4'h0; // @[Lookup.scala 33:37]
  wire [4:0] _T_543 = _T_269 ? 5'h1e : {{1'd0}, _T_542}; // @[Lookup.scala 33:37]
  wire [4:0] _T_544 = _T_267 ? 5'h1b : _T_543; // @[Lookup.scala 33:37]
  wire [6:0] _T_545 = _T_265 ? 7'h7b : {{2'd0}, _T_544}; // @[Lookup.scala 33:37]
  wire [6:0] _T_546 = _T_263 ? 7'h2 : _T_545; // @[Lookup.scala 33:37]
  wire [6:0] _T_547 = _T_261 ? 7'h21 : _T_546; // @[Lookup.scala 33:37]
  wire [6:0] _T_548 = _T_259 ? 7'h19 : _T_547; // @[Lookup.scala 33:37]
  wire [6:0] _T_549 = _T_257 ? 7'h11 : _T_548; // @[Lookup.scala 33:37]
  wire [6:0] _T_550 = _T_255 ? 7'h9 : _T_549; // @[Lookup.scala 33:37]
  wire [6:0] _T_551 = _T_253 ? 7'h1 : _T_550; // @[Lookup.scala 33:37]
  wire [6:0] _T_552 = _T_251 ? 7'h4 : _T_551; // @[Lookup.scala 33:37]
  wire [6:0] _T_553 = _T_249 ? 7'h0 : _T_552; // @[Lookup.scala 33:37]
  wire [6:0] _T_554 = _T_247 ? 7'h1 : _T_553; // @[Lookup.scala 33:37]
  wire [6:0] _T_555 = _T_245 ? 7'h7 : _T_554; // @[Lookup.scala 33:37]
  wire [6:0] _T_556 = _T_243 ? 7'h6 : _T_555; // @[Lookup.scala 33:37]
  wire [6:0] _T_557 = _T_241 ? 7'h5 : _T_556; // @[Lookup.scala 33:37]
  wire [6:0] _T_558 = _T_239 ? 7'h3 : _T_557; // @[Lookup.scala 33:37]
  wire [6:0] _T_559 = _T_237 ? 7'h2 : _T_558; // @[Lookup.scala 33:37]
  wire [6:0] _T_560 = _T_235 ? 7'h1 : _T_559; // @[Lookup.scala 33:37]
  wire [6:0] _T_561 = _T_233 ? 7'h32 : _T_560; // @[Lookup.scala 33:37]
  wire [6:0] _T_562 = _T_231 ? 7'h31 : _T_561; // @[Lookup.scala 33:37]
  wire [6:0] _T_563 = _T_229 ? 7'h30 : _T_562; // @[Lookup.scala 33:37]
  wire [6:0] _T_564 = _T_227 ? 7'h37 : _T_563; // @[Lookup.scala 33:37]
  wire [6:0] _T_565 = _T_225 ? 7'h26 : _T_564; // @[Lookup.scala 33:37]
  wire [6:0] _T_566 = _T_223 ? 7'h25 : _T_565; // @[Lookup.scala 33:37]
  wire [6:0] _T_567 = _T_221 ? 7'h24 : _T_566; // @[Lookup.scala 33:37]
  wire [6:0] _T_568 = _T_219 ? 7'h63 : _T_567; // @[Lookup.scala 33:37]
  wire [6:0] _T_569 = _T_217 ? 7'h22 : _T_568; // @[Lookup.scala 33:37]
  wire [6:0] _T_570 = _T_215 ? 7'h21 : _T_569; // @[Lookup.scala 33:37]
  wire [6:0] _T_571 = _T_213 ? 7'h21 : _T_570; // @[Lookup.scala 33:37]
  wire [6:0] _T_572 = _T_211 ? 7'h20 : _T_571; // @[Lookup.scala 33:37]
  wire [6:0] _T_573 = _T_209 ? 7'h20 : _T_572; // @[Lookup.scala 33:37]
  wire [6:0] _T_574 = _T_207 ? 7'h2 : _T_573; // @[Lookup.scala 33:37]
  wire [6:0] _T_575 = _T_205 ? 7'h0 : _T_574; // @[Lookup.scala 33:37]
  wire [6:0] _T_576 = _T_203 ? 7'h40 : _T_575; // @[Lookup.scala 33:37]
  wire [6:0] _T_577 = _T_201 ? 7'h0 : _T_576; // @[Lookup.scala 33:37]
  wire [6:0] _T_578 = _T_199 ? 7'h0 : _T_577; // @[Lookup.scala 33:37]
  wire [6:0] _T_579 = _T_197 ? 7'h0 : _T_578; // @[Lookup.scala 33:37]
  wire [6:0] _T_580 = _T_195 ? 7'h0 : _T_579; // @[Lookup.scala 33:37]
  wire [6:0] _T_581 = _T_193 ? 7'hb : _T_580; // @[Lookup.scala 33:37]
  wire [6:0] _T_582 = _T_191 ? 7'ha : _T_581; // @[Lookup.scala 33:37]
  wire [6:0] _T_583 = _T_189 ? 7'h40 : _T_582; // @[Lookup.scala 33:37]
  wire [6:0] _T_584 = _T_187 ? 7'h5a : _T_583; // @[Lookup.scala 33:37]
  wire [6:0] _T_585 = _T_185 ? 7'h0 : _T_584; // @[Lookup.scala 33:37]
  wire [6:0] _T_586 = _T_183 ? 7'h40 : _T_585; // @[Lookup.scala 33:37]
  wire [6:0] _T_587 = _T_181 ? 7'h5a : _T_586; // @[Lookup.scala 33:37]
  wire [6:0] _T_588 = _T_179 ? 7'h3 : _T_587; // @[Lookup.scala 33:37]
  wire [6:0] _T_589 = _T_177 ? 7'h2 : _T_588; // @[Lookup.scala 33:37]
  wire [6:0] _T_590 = _T_175 ? 7'h1 : _T_589; // @[Lookup.scala 33:37]
  wire [6:0] _T_591 = _T_173 ? 7'h11 : _T_590; // @[Lookup.scala 33:37]
  wire [6:0] _T_592 = _T_171 ? 7'h10 : _T_591; // @[Lookup.scala 33:37]
  wire [6:0] _T_593 = _T_169 ? 7'h58 : _T_592; // @[Lookup.scala 33:37]
  wire [6:0] _T_594 = _T_167 ? 7'h60 : _T_593; // @[Lookup.scala 33:37]
  wire [6:0] _T_595 = _T_165 ? 7'h28 : _T_594; // @[Lookup.scala 33:37]
  wire [6:0] _T_596 = _T_163 ? 7'h7 : _T_595; // @[Lookup.scala 33:37]
  wire [6:0] _T_597 = _T_161 ? 7'h6 : _T_596; // @[Lookup.scala 33:37]
  wire [6:0] _T_598 = _T_159 ? 7'h4 : _T_597; // @[Lookup.scala 33:37]
  wire [6:0] _T_599 = _T_157 ? 7'h8 : _T_598; // @[Lookup.scala 33:37]
  wire [6:0] _T_600 = _T_155 ? 7'h7 : _T_599; // @[Lookup.scala 33:37]
  wire [6:0] _T_601 = _T_153 ? 7'hd : _T_600; // @[Lookup.scala 33:37]
  wire [6:0] _T_602 = _T_151 ? 7'h5 : _T_601; // @[Lookup.scala 33:37]
  wire [6:0] _T_603 = _T_149 ? 7'h40 : _T_602; // @[Lookup.scala 33:37]
  wire [6:0] _T_604 = _T_147 ? 7'h40 : _T_603; // @[Lookup.scala 33:37]
  wire [6:0] _T_605 = _T_145 ? 7'h40 : _T_604; // @[Lookup.scala 33:37]
  wire [6:0] _T_606 = _T_143 ? 7'h60 : _T_605; // @[Lookup.scala 33:37]
  wire [6:0] _T_607 = _T_141 ? 7'h40 : _T_606; // @[Lookup.scala 33:37]
  wire [6:0] _T_608 = _T_139 ? 7'h40 : _T_607; // @[Lookup.scala 33:37]
  wire [6:0] _T_609 = _T_137 ? 7'hb : _T_608; // @[Lookup.scala 33:37]
  wire [6:0] _T_610 = _T_135 ? 7'ha : _T_609; // @[Lookup.scala 33:37]
  wire [6:0] _T_611 = _T_133 ? 7'h3 : _T_610; // @[Lookup.scala 33:37]
  wire [6:0] _T_612 = _T_131 ? 7'h2 : _T_611; // @[Lookup.scala 33:37]
  wire [6:0] _T_613 = _T_129 ? 7'h40 : _T_612; // @[Lookup.scala 33:37]
  wire [6:0] _T_614 = _T_127 ? 7'h0 : _T_613; // @[Lookup.scala 33:37]
  wire [6:0] _T_615 = _T_125 ? 7'hf : _T_614; // @[Lookup.scala 33:37]
  wire [6:0] _T_616 = _T_123 ? 7'he : _T_615; // @[Lookup.scala 33:37]
  wire [6:0] _T_617 = _T_121 ? 7'hd : _T_616; // @[Lookup.scala 33:37]
  wire [6:0] _T_618 = _T_119 ? 7'hc : _T_617; // @[Lookup.scala 33:37]
  wire [6:0] _T_619 = _T_117 ? 7'h8 : _T_618; // @[Lookup.scala 33:37]
  wire [6:0] _T_620 = _T_115 ? 7'h7 : _T_619; // @[Lookup.scala 33:37]
  wire [6:0] _T_621 = _T_113 ? 7'h6 : _T_620; // @[Lookup.scala 33:37]
  wire [6:0] _T_622 = _T_111 ? 7'h5 : _T_621; // @[Lookup.scala 33:37]
  wire [6:0] _T_623 = _T_109 ? 7'h4 : _T_622; // @[Lookup.scala 33:37]
  wire [6:0] _T_624 = _T_107 ? 7'h3 : _T_623; // @[Lookup.scala 33:37]
  wire [6:0] _T_625 = _T_105 ? 7'h2 : _T_624; // @[Lookup.scala 33:37]
  wire [6:0] _T_626 = _T_103 ? 7'h1 : _T_625; // @[Lookup.scala 33:37]
  wire [6:0] _T_627 = _T_101 ? 7'h0 : _T_626; // @[Lookup.scala 33:37]
  wire [6:0] _T_628 = _T_99 ? 7'h2 : _T_627; // @[Lookup.scala 33:37]
  wire [6:0] _T_629 = _T_97 ? 7'hb : _T_628; // @[Lookup.scala 33:37]
  wire [6:0] _T_630 = _T_95 ? 7'h3 : _T_629; // @[Lookup.scala 33:37]
  wire [6:0] _T_631 = _T_93 ? 7'h6 : _T_630; // @[Lookup.scala 33:37]
  wire [6:0] _T_632 = _T_91 ? 7'h28 : _T_631; // @[Lookup.scala 33:37]
  wire [6:0] _T_633 = _T_89 ? 7'h60 : _T_632; // @[Lookup.scala 33:37]
  wire [6:0] _T_634 = _T_87 ? 7'h2d : _T_633; // @[Lookup.scala 33:37]
  wire [6:0] _T_635 = _T_85 ? 7'h25 : _T_634; // @[Lookup.scala 33:37]
  wire [6:0] _T_636 = _T_83 ? 7'h21 : _T_635; // @[Lookup.scala 33:37]
  wire [6:0] _T_637 = _T_81 ? 7'h2d : _T_636; // @[Lookup.scala 33:37]
  wire [6:0] _T_638 = _T_79 ? 7'h25 : _T_637; // @[Lookup.scala 33:37]
  wire [6:0] _T_639 = _T_77 ? 7'h21 : _T_638; // @[Lookup.scala 33:37]
  wire [6:0] _T_640 = _T_75 ? 7'h60 : _T_639; // @[Lookup.scala 33:37]
  wire [6:0] _T_641 = _T_73 ? 7'ha : _T_640; // @[Lookup.scala 33:37]
  wire [6:0] _T_642 = _T_71 ? 7'h9 : _T_641; // @[Lookup.scala 33:37]
  wire [6:0] _T_643 = _T_69 ? 7'h8 : _T_642; // @[Lookup.scala 33:37]
  wire [6:0] _T_644 = _T_67 ? 7'h5 : _T_643; // @[Lookup.scala 33:37]
  wire [6:0] _T_645 = _T_65 ? 7'h4 : _T_644; // @[Lookup.scala 33:37]
  wire [6:0] _T_646 = _T_63 ? 7'h2 : _T_645; // @[Lookup.scala 33:37]
  wire [6:0] _T_647 = _T_61 ? 7'h1 : _T_646; // @[Lookup.scala 33:37]
  wire [6:0] _T_648 = _T_59 ? 7'h0 : _T_647; // @[Lookup.scala 33:37]
  wire [6:0] _T_649 = _T_57 ? 7'h17 : _T_648; // @[Lookup.scala 33:37]
  wire [6:0] _T_650 = _T_55 ? 7'h16 : _T_649; // @[Lookup.scala 33:37]
  wire [6:0] _T_651 = _T_53 ? 7'h15 : _T_650; // @[Lookup.scala 33:37]
  wire [6:0] _T_652 = _T_51 ? 7'h14 : _T_651; // @[Lookup.scala 33:37]
  wire [6:0] _T_653 = _T_49 ? 7'h11 : _T_652; // @[Lookup.scala 33:37]
  wire [6:0] _T_654 = _T_47 ? 7'h10 : _T_653; // @[Lookup.scala 33:37]
  wire [6:0] _T_655 = _T_45 ? 7'h5a : _T_654; // @[Lookup.scala 33:37]
  wire [6:0] _T_656 = _T_43 ? 7'h58 : _T_655; // @[Lookup.scala 33:37]
  wire [6:0] _T_657 = _T_41 ? 7'h40 : _T_656; // @[Lookup.scala 33:37]
  wire [6:0] _T_658 = _T_39 ? 7'h40 : _T_657; // @[Lookup.scala 33:37]
  wire [6:0] _T_659 = _T_37 ? 7'hd : _T_658; // @[Lookup.scala 33:37]
  wire [6:0] _T_660 = _T_35 ? 7'h8 : _T_659; // @[Lookup.scala 33:37]
  wire [6:0] _T_661 = _T_33 ? 7'h7 : _T_660; // @[Lookup.scala 33:37]
  wire [6:0] _T_662 = _T_31 ? 7'h6 : _T_661; // @[Lookup.scala 33:37]
  wire [6:0] _T_663 = _T_29 ? 7'h5 : _T_662; // @[Lookup.scala 33:37]
  wire [6:0] _T_664 = _T_27 ? 7'h4 : _T_663; // @[Lookup.scala 33:37]
  wire [6:0] _T_665 = _T_25 ? 7'h3 : _T_664; // @[Lookup.scala 33:37]
  wire [6:0] _T_666 = _T_23 ? 7'h2 : _T_665; // @[Lookup.scala 33:37]
  wire [6:0] _T_667 = _T_21 ? 7'h1 : _T_666; // @[Lookup.scala 33:37]
  wire [6:0] _T_668 = _T_19 ? 7'h40 : _T_667; // @[Lookup.scala 33:37]
  wire [6:0] _T_669 = _T_17 ? 7'hd : _T_668; // @[Lookup.scala 33:37]
  wire [6:0] _T_670 = _T_15 ? 7'h7 : _T_669; // @[Lookup.scala 33:37]
  wire [6:0] _T_671 = _T_13 ? 7'h6 : _T_670; // @[Lookup.scala 33:37]
  wire [6:0] _T_672 = _T_11 ? 7'h5 : _T_671; // @[Lookup.scala 33:37]
  wire [6:0] _T_673 = _T_9 ? 7'h4 : _T_672; // @[Lookup.scala 33:37]
  wire [6:0] _T_674 = _T_7 ? 7'h3 : _T_673; // @[Lookup.scala 33:37]
  wire [6:0] _T_675 = _T_5 ? 7'h2 : _T_674; // @[Lookup.scala 33:37]
  wire [6:0] _T_676 = _T_3 ? 7'h1 : _T_675; // @[Lookup.scala 33:37]
  wire [6:0] decodeList_2 = _T_1 ? 7'h40 : _T_676; // @[Lookup.scala 33:37]
  wire  hasIntr = |intrVecIDU; // @[IDU.scala 180:22]
  wire  _T_677 = hasIntr | io_in_bits_exceptionVec_12; // @[IDU.scala 36:84]
  wire  _T_678 = _T_677 | io_out_bits_cf_exceptionVec_1; // @[IDU.scala 36:127]
  wire [4:0] instrType = _T_678 ? 5'h0 : decodeList_0; // @[IDU.scala 36:75]
  wire [2:0] fuType = _T_678 ? 3'h3 : decodeList_1; // @[IDU.scala 36:75]
  wire [6:0] fuOpType = _T_678 ? 7'h0 : decodeList_2; // @[IDU.scala 36:75]
  wire  isRVC = io_in_bits_instr[1:0] != 2'h3; // @[IDU.scala 38:45]
  wire [4:0] _T_750 = _T_193 ? 5'h3 : 5'h10; // @[Lookup.scala 33:37]
  wire [4:0] _T_751 = _T_191 ? 5'h2 : _T_750; // @[Lookup.scala 33:37]
  wire [4:0] _T_752 = _T_189 ? 5'h10 : _T_751; // @[Lookup.scala 33:37]
  wire [4:0] _T_753 = _T_187 ? 5'h10 : _T_752; // @[Lookup.scala 33:37]
  wire [4:0] _T_754 = _T_185 ? 5'hf : _T_753; // @[Lookup.scala 33:37]
  wire [4:0] _T_755 = _T_183 ? 5'h10 : _T_754; // @[Lookup.scala 33:37]
  wire [4:0] _T_756 = _T_181 ? 5'h10 : _T_755; // @[Lookup.scala 33:37]
  wire [4:0] _T_757 = _T_179 ? 5'h1 : _T_756; // @[Lookup.scala 33:37]
  wire [4:0] _T_758 = _T_177 ? 5'h0 : _T_757; // @[Lookup.scala 33:37]
  wire [4:0] _T_759 = _T_175 ? 5'ha : _T_758; // @[Lookup.scala 33:37]
  wire [4:0] _T_760 = _T_173 ? 5'h9 : _T_759; // @[Lookup.scala 33:37]
  wire [4:0] _T_761 = _T_171 ? 5'h9 : _T_760; // @[Lookup.scala 33:37]
  wire [4:0] _T_762 = _T_169 ? 5'h8 : _T_761; // @[Lookup.scala 33:37]
  wire [4:0] _T_763 = _T_167 ? 5'h10 : _T_762; // @[Lookup.scala 33:37]
  wire [4:0] _T_764 = _T_165 ? 5'h10 : _T_763; // @[Lookup.scala 33:37]
  wire [4:0] _T_765 = _T_163 ? 5'h10 : _T_764; // @[Lookup.scala 33:37]
  wire [4:0] _T_766 = _T_161 ? 5'h10 : _T_765; // @[Lookup.scala 33:37]
  wire [4:0] _T_767 = _T_159 ? 5'h10 : _T_766; // @[Lookup.scala 33:37]
  wire [4:0] _T_768 = _T_157 ? 5'h10 : _T_767; // @[Lookup.scala 33:37]
  wire [4:0] _T_769 = _T_155 ? 5'ha : _T_768; // @[Lookup.scala 33:37]
  wire [4:0] _T_770 = _T_153 ? 5'ha : _T_769; // @[Lookup.scala 33:37]
  wire [4:0] _T_771 = _T_151 ? 5'ha : _T_770; // @[Lookup.scala 33:37]
  wire [4:0] _T_772 = _T_149 ? 5'hb : _T_771; // @[Lookup.scala 33:37]
  wire [4:0] _T_773 = _T_147 ? 5'hd : _T_772; // @[Lookup.scala 33:37]
  wire [4:0] _T_774 = _T_145 ? 5'ha : _T_773; // @[Lookup.scala 33:37]
  wire [4:0] _T_775 = _T_143 ? 5'hc : _T_774; // @[Lookup.scala 33:37]
  wire [4:0] _T_776 = _T_141 ? 5'hc : _T_775; // @[Lookup.scala 33:37]
  wire [4:0] _T_777 = _T_139 ? 5'h10 : _T_776; // @[Lookup.scala 33:37]
  wire [4:0] _T_778 = _T_137 ? 5'h5 : _T_777; // @[Lookup.scala 33:37]
  wire [4:0] _T_779 = _T_135 ? 5'h4 : _T_778; // @[Lookup.scala 33:37]
  wire [4:0] _T_780 = _T_133 ? 5'h7 : _T_779; // @[Lookup.scala 33:37]
  wire [4:0] _T_781 = _T_131 ? 5'h6 : _T_780; // @[Lookup.scala 33:37]
  wire [4:0] rvcImmType = _T_129 ? 5'he : _T_781; // @[Lookup.scala 33:37]
  wire [3:0] _T_782 = _T_193 ? 4'h9 : 4'h0; // @[Lookup.scala 33:37]
  wire [3:0] _T_783 = _T_191 ? 4'h9 : _T_782; // @[Lookup.scala 33:37]
  wire [3:0] _T_784 = _T_189 ? 4'h2 : _T_783; // @[Lookup.scala 33:37]
  wire [3:0] _T_785 = _T_187 ? 4'h4 : _T_784; // @[Lookup.scala 33:37]
  wire [3:0] _T_786 = _T_185 ? 4'h0 : _T_785; // @[Lookup.scala 33:37]
  wire [3:0] _T_787 = _T_183 ? 4'h5 : _T_786; // @[Lookup.scala 33:37]
  wire [3:0] _T_788 = _T_181 ? 4'h4 : _T_787; // @[Lookup.scala 33:37]
  wire [3:0] _T_789 = _T_179 ? 4'h9 : _T_788; // @[Lookup.scala 33:37]
  wire [3:0] _T_790 = _T_177 ? 4'h9 : _T_789; // @[Lookup.scala 33:37]
  wire [3:0] _T_791 = _T_175 ? 4'h2 : _T_790; // @[Lookup.scala 33:37]
  wire [3:0] _T_792 = _T_173 ? 4'h6 : _T_791; // @[Lookup.scala 33:37]
  wire [3:0] _T_793 = _T_171 ? 4'h6 : _T_792; // @[Lookup.scala 33:37]
  wire [3:0] _T_794 = _T_169 ? 4'h0 : _T_793; // @[Lookup.scala 33:37]
  wire [3:0] _T_795 = _T_167 ? 4'h6 : _T_794; // @[Lookup.scala 33:37]
  wire [3:0] _T_796 = _T_165 ? 4'h6 : _T_795; // @[Lookup.scala 33:37]
  wire [3:0] _T_797 = _T_163 ? 4'h6 : _T_796; // @[Lookup.scala 33:37]
  wire [3:0] _T_798 = _T_161 ? 4'h6 : _T_797; // @[Lookup.scala 33:37]
  wire [3:0] _T_799 = _T_159 ? 4'h6 : _T_798; // @[Lookup.scala 33:37]
  wire [3:0] _T_800 = _T_157 ? 4'h6 : _T_799; // @[Lookup.scala 33:37]
  wire [3:0] _T_801 = _T_155 ? 4'h6 : _T_800; // @[Lookup.scala 33:37]
  wire [3:0] _T_802 = _T_153 ? 4'h6 : _T_801; // @[Lookup.scala 33:37]
  wire [3:0] _T_803 = _T_151 ? 4'h6 : _T_802; // @[Lookup.scala 33:37]
  wire [3:0] _T_804 = _T_149 ? 4'h0 : _T_803; // @[Lookup.scala 33:37]
  wire [3:0] _T_805 = _T_147 ? 4'h9 : _T_804; // @[Lookup.scala 33:37]
  wire [3:0] _T_806 = _T_145 ? 4'h0 : _T_805; // @[Lookup.scala 33:37]
  wire [3:0] _T_807 = _T_143 ? 4'h2 : _T_806; // @[Lookup.scala 33:37]
  wire [3:0] _T_808 = _T_141 ? 4'h2 : _T_807; // @[Lookup.scala 33:37]
  wire [3:0] _T_809 = _T_139 ? 4'h0 : _T_808; // @[Lookup.scala 33:37]
  wire [3:0] _T_810 = _T_137 ? 4'h6 : _T_809; // @[Lookup.scala 33:37]
  wire [3:0] _T_811 = _T_135 ? 4'h6 : _T_810; // @[Lookup.scala 33:37]
  wire [3:0] _T_812 = _T_133 ? 4'h6 : _T_811; // @[Lookup.scala 33:37]
  wire [3:0] _T_813 = _T_131 ? 4'h6 : _T_812; // @[Lookup.scala 33:37]
  wire [3:0] rvcSrc1Type = _T_129 ? 4'h9 : _T_813; // @[Lookup.scala 33:37]
  wire [2:0] _T_814 = _T_193 ? 3'h5 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _T_815 = _T_191 ? 3'h5 : _T_814; // @[Lookup.scala 33:37]
  wire [2:0] _T_816 = _T_189 ? 3'h5 : _T_815; // @[Lookup.scala 33:37]
  wire [2:0] _T_817 = _T_187 ? 3'h0 : _T_816; // @[Lookup.scala 33:37]
  wire [2:0] _T_818 = _T_185 ? 3'h0 : _T_817; // @[Lookup.scala 33:37]
  wire [2:0] _T_819 = _T_183 ? 3'h0 : _T_818; // @[Lookup.scala 33:37]
  wire [2:0] _T_820 = _T_181 ? 3'h0 : _T_819; // @[Lookup.scala 33:37]
  wire [2:0] _T_821 = _T_179 ? 3'h0 : _T_820; // @[Lookup.scala 33:37]
  wire [2:0] _T_822 = _T_177 ? 3'h0 : _T_821; // @[Lookup.scala 33:37]
  wire [2:0] _T_823 = _T_175 ? 3'h0 : _T_822; // @[Lookup.scala 33:37]
  wire [2:0] _T_824 = _T_173 ? 3'h0 : _T_823; // @[Lookup.scala 33:37]
  wire [2:0] _T_825 = _T_171 ? 3'h0 : _T_824; // @[Lookup.scala 33:37]
  wire [2:0] _T_826 = _T_169 ? 3'h0 : _T_825; // @[Lookup.scala 33:37]
  wire [2:0] _T_827 = _T_167 ? 3'h7 : _T_826; // @[Lookup.scala 33:37]
  wire [2:0] _T_828 = _T_165 ? 3'h7 : _T_827; // @[Lookup.scala 33:37]
  wire [2:0] _T_829 = _T_163 ? 3'h7 : _T_828; // @[Lookup.scala 33:37]
  wire [2:0] _T_830 = _T_161 ? 3'h7 : _T_829; // @[Lookup.scala 33:37]
  wire [2:0] _T_831 = _T_159 ? 3'h7 : _T_830; // @[Lookup.scala 33:37]
  wire [2:0] _T_832 = _T_157 ? 3'h7 : _T_831; // @[Lookup.scala 33:37]
  wire [2:0] _T_833 = _T_155 ? 3'h0 : _T_832; // @[Lookup.scala 33:37]
  wire [2:0] _T_834 = _T_153 ? 3'h0 : _T_833; // @[Lookup.scala 33:37]
  wire [2:0] _T_835 = _T_151 ? 3'h0 : _T_834; // @[Lookup.scala 33:37]
  wire [2:0] _T_836 = _T_149 ? 3'h0 : _T_835; // @[Lookup.scala 33:37]
  wire [2:0] _T_837 = _T_147 ? 3'h0 : _T_836; // @[Lookup.scala 33:37]
  wire [2:0] _T_838 = _T_145 ? 3'h0 : _T_837; // @[Lookup.scala 33:37]
  wire [2:0] _T_839 = _T_143 ? 3'h0 : _T_838; // @[Lookup.scala 33:37]
  wire [2:0] _T_840 = _T_141 ? 3'h0 : _T_839; // @[Lookup.scala 33:37]
  wire [2:0] _T_841 = _T_139 ? 3'h0 : _T_840; // @[Lookup.scala 33:37]
  wire [2:0] _T_842 = _T_137 ? 3'h7 : _T_841; // @[Lookup.scala 33:37]
  wire [2:0] _T_843 = _T_135 ? 3'h7 : _T_842; // @[Lookup.scala 33:37]
  wire [2:0] _T_844 = _T_133 ? 3'h0 : _T_843; // @[Lookup.scala 33:37]
  wire [2:0] _T_845 = _T_131 ? 3'h0 : _T_844; // @[Lookup.scala 33:37]
  wire [2:0] rvcSrc2Type = _T_129 ? 3'h0 : _T_845; // @[Lookup.scala 33:37]
  wire [1:0] _T_848 = _T_189 ? 2'h2 : 2'h0; // @[Lookup.scala 33:37]
  wire [3:0] _T_849 = _T_187 ? 4'h8 : {{2'd0}, _T_848}; // @[Lookup.scala 33:37]
  wire [3:0] _T_850 = _T_185 ? 4'h0 : _T_849; // @[Lookup.scala 33:37]
  wire [3:0] _T_851 = _T_183 ? 4'h2 : _T_850; // @[Lookup.scala 33:37]
  wire [3:0] _T_852 = _T_181 ? 4'h0 : _T_851; // @[Lookup.scala 33:37]
  wire [3:0] _T_853 = _T_179 ? 4'h2 : _T_852; // @[Lookup.scala 33:37]
  wire [3:0] _T_854 = _T_177 ? 4'h2 : _T_853; // @[Lookup.scala 33:37]
  wire [3:0] _T_855 = _T_175 ? 4'h2 : _T_854; // @[Lookup.scala 33:37]
  wire [3:0] _T_856 = _T_173 ? 4'h0 : _T_855; // @[Lookup.scala 33:37]
  wire [3:0] _T_857 = _T_171 ? 4'h0 : _T_856; // @[Lookup.scala 33:37]
  wire [3:0] _T_858 = _T_169 ? 4'h0 : _T_857; // @[Lookup.scala 33:37]
  wire [3:0] _T_859 = _T_167 ? 4'h6 : _T_858; // @[Lookup.scala 33:37]
  wire [3:0] _T_860 = _T_165 ? 4'h6 : _T_859; // @[Lookup.scala 33:37]
  wire [3:0] _T_861 = _T_163 ? 4'h6 : _T_860; // @[Lookup.scala 33:37]
  wire [3:0] _T_862 = _T_161 ? 4'h6 : _T_861; // @[Lookup.scala 33:37]
  wire [3:0] _T_863 = _T_159 ? 4'h6 : _T_862; // @[Lookup.scala 33:37]
  wire [3:0] _T_864 = _T_157 ? 4'h6 : _T_863; // @[Lookup.scala 33:37]
  wire [3:0] _T_865 = _T_155 ? 4'h6 : _T_864; // @[Lookup.scala 33:37]
  wire [3:0] _T_866 = _T_153 ? 4'h6 : _T_865; // @[Lookup.scala 33:37]
  wire [3:0] _T_867 = _T_151 ? 4'h6 : _T_866; // @[Lookup.scala 33:37]
  wire [3:0] _T_868 = _T_149 ? 4'h2 : _T_867; // @[Lookup.scala 33:37]
  wire [3:0] _T_869 = _T_147 ? 4'h9 : _T_868; // @[Lookup.scala 33:37]
  wire [3:0] _T_870 = _T_145 ? 4'h2 : _T_869; // @[Lookup.scala 33:37]
  wire [3:0] _T_871 = _T_143 ? 4'h2 : _T_870; // @[Lookup.scala 33:37]
  wire [3:0] _T_872 = _T_141 ? 4'h2 : _T_871; // @[Lookup.scala 33:37]
  wire [3:0] _T_873 = _T_139 ? 4'h0 : _T_872; // @[Lookup.scala 33:37]
  wire [3:0] _T_874 = _T_137 ? 4'h0 : _T_873; // @[Lookup.scala 33:37]
  wire [3:0] _T_875 = _T_135 ? 4'h0 : _T_874; // @[Lookup.scala 33:37]
  wire [3:0] _T_876 = _T_133 ? 4'h7 : _T_875; // @[Lookup.scala 33:37]
  wire [3:0] _T_877 = _T_131 ? 4'h7 : _T_876; // @[Lookup.scala 33:37]
  wire [3:0] rvcDestType = _T_129 ? 4'h7 : _T_877; // @[Lookup.scala 33:37]
  wire  _T_878 = 5'h4 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_880 = 5'h2 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_881 = 5'hf == instrType; // @[LookupTree.scala 24:34]
  wire  _T_882 = 5'h1 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_883 = 5'h6 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_884 = 5'h7 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_885 = 5'h0 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_886 = 5'h10 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_887 = 5'h15 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_888 = 5'h16 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_889 = 5'h17 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_907 = _T_883 | _T_884; // @[Mux.scala 27:72]
  wire  _T_908 = _T_907 | _T_885; // @[Mux.scala 27:72]
  wire  src1Type = _T_908 | _T_889; // @[Mux.scala 27:72]
  wire  _T_941 = _T_878 | _T_883; // @[Mux.scala 27:72]
  wire  _T_942 = _T_941 | _T_884; // @[Mux.scala 27:72]
  wire  _T_943 = _T_942 | _T_885; // @[Mux.scala 27:72]
  wire  _T_945 = _T_943 | _T_887; // @[Mux.scala 27:72]
  wire  src2Type = _T_945 | _T_889; // @[Mux.scala 27:72]
  wire [4:0] rs = io_in_bits_instr[19:15]; // @[IDU.scala 64:28]
  wire [4:0] rt = io_in_bits_instr[24:20]; // @[IDU.scala 64:43]
  wire [4:0] rd = io_in_bits_instr[11:7]; // @[IDU.scala 64:58]
  wire [4:0] rs2 = io_in_bits_instr[6:2]; // @[IDU.scala 68:24]
  wire  _T_949 = 3'h0 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_950 = 3'h1 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_951 = 3'h2 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_952 = 3'h3 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_953 = 3'h4 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_954 = 3'h5 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_955 = 3'h6 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_956 = 3'h7 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire [3:0] _T_957 = _T_949 ? 4'h8 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_958 = _T_950 ? 4'h9 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_959 = _T_951 ? 4'ha : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_960 = _T_952 ? 4'hb : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_961 = _T_953 ? 4'hc : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_962 = _T_954 ? 4'hd : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_963 = _T_955 ? 4'he : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_964 = _T_956 ? 4'hf : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_965 = _T_957 | _T_958; // @[Mux.scala 27:72]
  wire [3:0] _T_966 = _T_965 | _T_959; // @[Mux.scala 27:72]
  wire [3:0] _T_967 = _T_966 | _T_960; // @[Mux.scala 27:72]
  wire [3:0] _T_968 = _T_967 | _T_961; // @[Mux.scala 27:72]
  wire [3:0] _T_969 = _T_968 | _T_962; // @[Mux.scala 27:72]
  wire [3:0] _T_970 = _T_969 | _T_963; // @[Mux.scala 27:72]
  wire [3:0] rs1p = _T_970 | _T_964; // @[Mux.scala 27:72]
  wire  _T_973 = 3'h0 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_974 = 3'h1 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_975 = 3'h2 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_976 = 3'h3 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_977 = 3'h4 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_978 = 3'h5 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_979 = 3'h6 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_980 = 3'h7 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire [3:0] _T_981 = _T_973 ? 4'h8 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_982 = _T_974 ? 4'h9 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_983 = _T_975 ? 4'ha : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_984 = _T_976 ? 4'hb : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_985 = _T_977 ? 4'hc : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_986 = _T_978 ? 4'hd : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_987 = _T_979 ? 4'he : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_988 = _T_980 ? 4'hf : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_989 = _T_981 | _T_982; // @[Mux.scala 27:72]
  wire [3:0] _T_990 = _T_989 | _T_983; // @[Mux.scala 27:72]
  wire [3:0] _T_991 = _T_990 | _T_984; // @[Mux.scala 27:72]
  wire [3:0] _T_992 = _T_991 | _T_985; // @[Mux.scala 27:72]
  wire [3:0] _T_993 = _T_992 | _T_986; // @[Mux.scala 27:72]
  wire [3:0] _T_994 = _T_993 | _T_987; // @[Mux.scala 27:72]
  wire [3:0] rs2p = _T_994 | _T_988; // @[Mux.scala 27:72]
  wire [5:0] rvc_shamt = {io_in_bits_instr[12],rs2}; // @[Cat.scala 29:58]
  wire  _T_999 = 4'h3 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_1000 = 4'h1 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_1001 = 4'h2 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_1002 = 4'h4 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_1003 = 4'h5 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_1004 = 4'h6 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_1005 = 4'h7 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_1006 = 4'h8 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_1007 = 4'h9 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire [4:0] _T_1009 = _T_999 ? rs : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1010 = _T_1000 ? rt : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1011 = _T_1001 ? rd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1012 = _T_1002 ? rd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1013 = _T_1003 ? rs2 : 5'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_1014 = _T_1004 ? rs1p : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_1015 = _T_1005 ? rs2p : 4'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_1017 = _T_1007 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1019 = _T_1009 | _T_1010; // @[Mux.scala 27:72]
  wire [4:0] _T_1020 = _T_1019 | _T_1011; // @[Mux.scala 27:72]
  wire [4:0] _T_1021 = _T_1020 | _T_1012; // @[Mux.scala 27:72]
  wire [4:0] _T_1022 = _T_1021 | _T_1013; // @[Mux.scala 27:72]
  wire [4:0] _GEN_5 = {{1'd0}, _T_1014}; // @[Mux.scala 27:72]
  wire [4:0] _T_1023 = _T_1022 | _GEN_5; // @[Mux.scala 27:72]
  wire [4:0] _GEN_6 = {{1'd0}, _T_1015}; // @[Mux.scala 27:72]
  wire [4:0] _T_1024 = _T_1023 | _GEN_6; // @[Mux.scala 27:72]
  wire [4:0] _GEN_7 = {{4'd0}, _T_1006}; // @[Mux.scala 27:72]
  wire [4:0] _T_1025 = _T_1024 | _GEN_7; // @[Mux.scala 27:72]
  wire [4:0] _GEN_8 = {{3'd0}, _T_1017}; // @[Mux.scala 27:72]
  wire [4:0] rvc_src1 = _T_1025 | _GEN_8; // @[Mux.scala 27:72]
  wire  _T_1028 = 3'h3 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire  _T_1029 = 3'h1 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire  _T_1030 = 3'h2 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire  _T_1031 = 3'h4 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire  _T_1032 = 3'h5 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire  _T_1033 = 3'h6 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire  _T_1034 = 3'h7 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire [3:0] _GEN_9 = {{1'd0}, rvcSrc2Type}; // @[LookupTree.scala 24:34]
  wire  _T_1035 = 4'h8 == _GEN_9; // @[LookupTree.scala 24:34]
  wire  _T_1036 = 4'h9 == _GEN_9; // @[LookupTree.scala 24:34]
  wire [4:0] _T_1038 = _T_1028 ? rs : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1039 = _T_1029 ? rt : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1040 = _T_1030 ? rd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1041 = _T_1031 ? rd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1042 = _T_1032 ? rs2 : 5'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_1043 = _T_1033 ? rs1p : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_1044 = _T_1034 ? rs2p : 4'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_1046 = _T_1036 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1048 = _T_1038 | _T_1039; // @[Mux.scala 27:72]
  wire [4:0] _T_1049 = _T_1048 | _T_1040; // @[Mux.scala 27:72]
  wire [4:0] _T_1050 = _T_1049 | _T_1041; // @[Mux.scala 27:72]
  wire [4:0] _T_1051 = _T_1050 | _T_1042; // @[Mux.scala 27:72]
  wire [4:0] _GEN_11 = {{1'd0}, _T_1043}; // @[Mux.scala 27:72]
  wire [4:0] _T_1052 = _T_1051 | _GEN_11; // @[Mux.scala 27:72]
  wire [4:0] _GEN_12 = {{1'd0}, _T_1044}; // @[Mux.scala 27:72]
  wire [4:0] _T_1053 = _T_1052 | _GEN_12; // @[Mux.scala 27:72]
  wire [4:0] _GEN_13 = {{4'd0}, _T_1035}; // @[Mux.scala 27:72]
  wire [4:0] _T_1054 = _T_1053 | _GEN_13; // @[Mux.scala 27:72]
  wire [4:0] _GEN_14 = {{3'd0}, _T_1046}; // @[Mux.scala 27:72]
  wire [4:0] rvc_src2 = _T_1054 | _GEN_14; // @[Mux.scala 27:72]
  wire  _T_1057 = 4'h3 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_1058 = 4'h1 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_1059 = 4'h2 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_1060 = 4'h4 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_1061 = 4'h5 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_1062 = 4'h6 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_1063 = 4'h7 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_1064 = 4'h8 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_1065 = 4'h9 == rvcDestType; // @[LookupTree.scala 24:34]
  wire [4:0] _T_1067 = _T_1057 ? rs : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1068 = _T_1058 ? rt : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1069 = _T_1059 ? rd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1070 = _T_1060 ? rd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1071 = _T_1061 ? rs2 : 5'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_1072 = _T_1062 ? rs1p : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_1073 = _T_1063 ? rs2p : 4'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_1075 = _T_1065 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1077 = _T_1067 | _T_1068; // @[Mux.scala 27:72]
  wire [4:0] _T_1078 = _T_1077 | _T_1069; // @[Mux.scala 27:72]
  wire [4:0] _T_1079 = _T_1078 | _T_1070; // @[Mux.scala 27:72]
  wire [4:0] _T_1080 = _T_1079 | _T_1071; // @[Mux.scala 27:72]
  wire [4:0] _GEN_15 = {{1'd0}, _T_1072}; // @[Mux.scala 27:72]
  wire [4:0] _T_1081 = _T_1080 | _GEN_15; // @[Mux.scala 27:72]
  wire [4:0] _GEN_16 = {{1'd0}, _T_1073}; // @[Mux.scala 27:72]
  wire [4:0] _T_1082 = _T_1081 | _GEN_16; // @[Mux.scala 27:72]
  wire [4:0] _GEN_17 = {{4'd0}, _T_1064}; // @[Mux.scala 27:72]
  wire [4:0] _T_1083 = _T_1082 | _GEN_17; // @[Mux.scala 27:72]
  wire [4:0] _GEN_18 = {{3'd0}, _T_1075}; // @[Mux.scala 27:72]
  wire [4:0] rvc_dest = _T_1083 | _GEN_18; // @[Mux.scala 27:72]
  wire [4:0] rfSrc1 = isRVC ? rvc_src1 : rs; // @[IDU.scala 92:19]
  wire [4:0] rfSrc2 = isRVC ? rvc_src2 : rt; // @[IDU.scala 93:19]
  wire [4:0] rfDest = isRVC ? rvc_dest : rd; // @[IDU.scala 94:19]
  wire  _T_1087 = ~src2Type; // @[IDU.scala 98:43]
  wire [51:0] _T_1095 = io_in_bits_instr[31] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1096 = {_T_1095,io_in_bits_instr[31:20]}; // @[Cat.scala 29:58]
  wire [11:0] _T_1099 = {io_in_bits_instr[31:25],rd}; // @[Cat.scala 29:58]
  wire [51:0] _T_1102 = _T_1099[11] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1103 = {_T_1102,io_in_bits_instr[31:25],rd}; // @[Cat.scala 29:58]
  wire [12:0] _T_1118 = {io_in_bits_instr[31],io_in_bits_instr[7],io_in_bits_instr[30:25],io_in_bits_instr[11:8],1'h0}; // @[Cat.scala 29:58]
  wire [50:0] _T_1121 = _T_1118[12] ? 51'h7ffffffffffff : 51'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1122 = {_T_1121,io_in_bits_instr[31],io_in_bits_instr[7],io_in_bits_instr[30:25],io_in_bits_instr[11:8],1'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_1124 = {io_in_bits_instr[31:12],12'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_1127 = _T_1124[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1128 = {_T_1127,io_in_bits_instr[31:12],12'h0}; // @[Cat.scala 29:58]
  wire [20:0] _T_1136 = {io_in_bits_instr[31],io_in_bits_instr[19:12],io_in_bits_instr[20],io_in_bits_instr[30:21],1'h0}; // @[Cat.scala 29:58]
  wire [42:0] _T_1139 = _T_1136[20] ? 43'h7ffffffffff : 43'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1140 = {_T_1139,io_in_bits_instr[31],io_in_bits_instr[19:12],io_in_bits_instr[20],io_in_bits_instr[30:21],1'h0}; // @[Cat.scala 29:58]
  wire [63:0] _T_1142 = {57'h0,io_in_bits_instr[31:25]}; // @[Cat.scala 29:58]
  wire [63:0] _T_1144 = {52'h0,io_in_bits_instr[31:20]}; // @[Cat.scala 29:58]
  wire [63:0] _T_1148 = {52'h0,io_in_bits_instr[31:25],rd}; // @[Cat.scala 29:58]
  wire [63:0] _T_1151 = {35'h0,12'h0,io_in_bits_instr[31:15]}; // @[Cat.scala 29:58]
  wire [63:0] _T_1153 = {54'h0,io_in_bits_instr[24:15]}; // @[Cat.scala 29:58]
  wire  _T_1164 = 5'h1f == instrType; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1165 = _T_878 ? _T_1096 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1166 = _T_880 ? _T_1103 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1167 = _T_881 ? _T_1103 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1168 = _T_882 ? _T_1122 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1169 = _T_883 ? _T_1128 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1170 = _T_884 ? _T_1140 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1171 = _T_888 ? _T_1142 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1172 = _T_887 ? _T_1144 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1173 = _T_886 ? _T_1148 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1174 = _T_889 ? _T_1151 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1175 = _T_1164 ? _T_1153 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1176 = _T_1165 | _T_1166; // @[Mux.scala 27:72]
  wire [63:0] _T_1177 = _T_1176 | _T_1167; // @[Mux.scala 27:72]
  wire [63:0] _T_1178 = _T_1177 | _T_1168; // @[Mux.scala 27:72]
  wire [63:0] _T_1179 = _T_1178 | _T_1169; // @[Mux.scala 27:72]
  wire [63:0] _T_1180 = _T_1179 | _T_1170; // @[Mux.scala 27:72]
  wire [63:0] _T_1181 = _T_1180 | _T_1171; // @[Mux.scala 27:72]
  wire [63:0] _T_1182 = _T_1181 | _T_1172; // @[Mux.scala 27:72]
  wire [63:0] _T_1183 = _T_1182 | _T_1173; // @[Mux.scala 27:72]
  wire [63:0] _T_1184 = _T_1183 | _T_1174; // @[Mux.scala 27:72]
  wire [63:0] imm = _T_1184 | _T_1175; // @[Mux.scala 27:72]
  wire [63:0] _T_1192 = {56'h0,io_in_bits_instr[3:2],io_in_bits_instr[12],io_in_bits_instr[6:4],2'h0}; // @[Cat.scala 29:58]
  wire [63:0] _T_1199 = {55'h0,io_in_bits_instr[4:2],io_in_bits_instr[12],io_in_bits_instr[6:5],3'h0}; // @[Cat.scala 29:58]
  wire [63:0] _T_1204 = {56'h0,io_in_bits_instr[8:7],io_in_bits_instr[12:9],2'h0}; // @[Cat.scala 29:58]
  wire [63:0] _T_1209 = {55'h0,io_in_bits_instr[9:7],io_in_bits_instr[12:10],3'h0}; // @[Cat.scala 29:58]
  wire [63:0] _T_1216 = {57'h0,io_in_bits_instr[5],io_in_bits_instr[12:10],io_in_bits_instr[6],2'h0}; // @[Cat.scala 29:58]
  wire [63:0] _T_1221 = {56'h0,io_in_bits_instr[6:5],io_in_bits_instr[12:10],3'h0}; // @[Cat.scala 29:58]
  wire [11:0] _T_1249 = {io_in_bits_instr[12],io_in_bits_instr[8],io_in_bits_instr[10:9],io_in_bits_instr[6],io_in_bits_instr[7],io_in_bits_instr[2],io_in_bits_instr[11],io_in_bits_instr[5:3],1'h0}; // @[Cat.scala 29:58]
  wire [51:0] _T_1252 = _T_1249[11] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1253 = {_T_1252,io_in_bits_instr[12],io_in_bits_instr[8],io_in_bits_instr[10:9],io_in_bits_instr[6],io_in_bits_instr[7],io_in_bits_instr[2],io_in_bits_instr[11],io_in_bits_instr[5:3],1'h0}; // @[Cat.scala 29:58]
  wire [8:0] _T_1263 = {io_in_bits_instr[12],io_in_bits_instr[6:5],io_in_bits_instr[2],io_in_bits_instr[11:10],io_in_bits_instr[4:3],1'h0}; // @[Cat.scala 29:58]
  wire [54:0] _T_1266 = _T_1263[8] ? 55'h7fffffffffffff : 55'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1267 = {_T_1266,io_in_bits_instr[12],io_in_bits_instr[6:5],io_in_bits_instr[2],io_in_bits_instr[11:10],io_in_bits_instr[4:3],1'h0}; // @[Cat.scala 29:58]
  wire [57:0] _T_1273 = rvc_shamt[5] ? 58'h3ffffffffffffff : 58'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1274 = {_T_1273,io_in_bits_instr[12],rs2}; // @[Cat.scala 29:58]
  wire [17:0] _T_1278 = {io_in_bits_instr[12],rs2,12'h0}; // @[Cat.scala 29:58]
  wire [45:0] _T_1281 = _T_1278[17] ? 46'h3fffffffffff : 46'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1282 = {_T_1281,io_in_bits_instr[12],rs2,12'h0}; // @[Cat.scala 29:58]
  wire [9:0] _T_1299 = {io_in_bits_instr[12],io_in_bits_instr[4:3],io_in_bits_instr[5],io_in_bits_instr[2],io_in_bits_instr[6],4'h0}; // @[Cat.scala 29:58]
  wire [53:0] _T_1302 = _T_1299[9] ? 54'h3fffffffffffff : 54'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1303 = {_T_1302,io_in_bits_instr[12],io_in_bits_instr[4:3],io_in_bits_instr[5],io_in_bits_instr[2],io_in_bits_instr[6],4'h0}; // @[Cat.scala 29:58]
  wire [63:0] _T_1312 = {54'h0,io_in_bits_instr[10:7],io_in_bits_instr[12:11],io_in_bits_instr[5],io_in_bits_instr[6],2'h0}; // @[Cat.scala 29:58]
  wire  _T_1314 = 5'h0 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1315 = 5'h1 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1316 = 5'h2 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1317 = 5'h3 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1318 = 5'h4 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1319 = 5'h5 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1320 = 5'h6 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1321 = 5'h7 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1322 = 5'h8 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1323 = 5'h9 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1324 = 5'ha == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1325 = 5'hb == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1326 = 5'hc == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1327 = 5'hd == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1328 = 5'he == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1329 = 5'hf == rvcImmType; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1331 = _T_1314 ? _T_1192 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1332 = _T_1315 ? _T_1199 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1333 = _T_1316 ? _T_1204 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1334 = _T_1317 ? _T_1209 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1335 = _T_1318 ? _T_1216 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1336 = _T_1319 ? _T_1221 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1337 = _T_1320 ? _T_1216 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1338 = _T_1321 ? _T_1221 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1339 = _T_1322 ? _T_1253 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1340 = _T_1323 ? _T_1267 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1341 = _T_1324 ? _T_1274 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1342 = _T_1325 ? _T_1282 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1343 = _T_1326 ? _T_1274 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1344 = _T_1327 ? _T_1303 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1345 = _T_1328 ? _T_1312 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1346 = _T_1329 ? 64'h1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1348 = _T_1331 | _T_1332; // @[Mux.scala 27:72]
  wire [63:0] _T_1349 = _T_1348 | _T_1333; // @[Mux.scala 27:72]
  wire [63:0] _T_1350 = _T_1349 | _T_1334; // @[Mux.scala 27:72]
  wire [63:0] _T_1351 = _T_1350 | _T_1335; // @[Mux.scala 27:72]
  wire [63:0] _T_1352 = _T_1351 | _T_1336; // @[Mux.scala 27:72]
  wire [63:0] _T_1353 = _T_1352 | _T_1337; // @[Mux.scala 27:72]
  wire [63:0] _T_1354 = _T_1353 | _T_1338; // @[Mux.scala 27:72]
  wire [63:0] _T_1355 = _T_1354 | _T_1339; // @[Mux.scala 27:72]
  wire [63:0] _T_1356 = _T_1355 | _T_1340; // @[Mux.scala 27:72]
  wire [63:0] _T_1357 = _T_1356 | _T_1341; // @[Mux.scala 27:72]
  wire [63:0] _T_1358 = _T_1357 | _T_1342; // @[Mux.scala 27:72]
  wire [63:0] _T_1359 = _T_1358 | _T_1343; // @[Mux.scala 27:72]
  wire [63:0] _T_1360 = _T_1359 | _T_1344; // @[Mux.scala 27:72]
  wire [63:0] _T_1361 = _T_1360 | _T_1345; // @[Mux.scala 27:72]
  wire [63:0] immrvc = _T_1361 | _T_1346; // @[Mux.scala 27:72]
  wire  _T_1364 = fuType == 3'h0; // @[IDU.scala 140:16]
  wire  _T_1365 = rfDest == 5'h1; // @[IDU.scala 141:34]
  wire  _T_1366 = rfDest == 5'h5; // @[IDU.scala 141:49]
  wire  _T_1367 = _T_1365 | _T_1366; // @[IDU.scala 141:42]
  wire  _T_1368 = fuOpType == 7'h58; // @[IDU.scala 142:38]
  wire  _T_1369 = _T_1367 & _T_1368; // @[IDU.scala 142:26]
  wire [6:0] _GEN_0 = _T_1369 ? 7'h5c : fuOpType; // @[IDU.scala 142:57]
  wire  _T_1370 = fuOpType == 7'h5a; // @[IDU.scala 143:20]
  wire  _T_1371 = rfSrc1 == 5'h1; // @[IDU.scala 141:34]
  wire  _T_1372 = rfSrc1 == 5'h5; // @[IDU.scala 141:49]
  wire  _T_1373 = _T_1371 | _T_1372; // @[IDU.scala 141:42]
  wire [6:0] _GEN_1 = _T_1373 ? 7'h5e : _GEN_0; // @[IDU.scala 144:29]
  wire [6:0] _GEN_2 = _T_1367 ? 7'h5c : _GEN_1; // @[IDU.scala 145:29]
  wire [6:0] _GEN_3 = _T_1370 ? _GEN_2 : _GEN_0; // @[IDU.scala 143:40]
  wire  _T_1378 = io_in_bits_instr[6:0] == 7'h37; // @[IDU.scala 149:47]
  wire  _T_1379 = _T_1378 ? 1'h0 : src1Type; // @[IDU.scala 149:35]
  wire  _T_1390 = ~io_in_valid; // @[IDU.scala 170:18]
  wire  _T_1391 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_1392 = ~hasIntr; // @[IDU.scala 170:51]
  wire  _T_1393 = _T_1391 & _T_1392; // @[IDU.scala 170:48]
  reg [63:0] _T_1396; // @[GTimer.scala 24:20]
  wire [63:0] _T_1398 = _T_1396 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_1400 = _T_1391 & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  wire  _T_1402 = ~reset; // @[Debug.scala 56:24]
  wire  _T_1418 = instrType == 5'h0; // @[IDU.scala 186:59]
  wire  _T_1420 = _T_1418 & _T_1392; // @[IDU.scala 186:70]
  wire  _T_1423 = |io_in_bits_pc[38:32]; // @[IDU.scala 189:94]
  wire  _T_1424 = ~DTLBENABLE; // @[IDU.scala 189:101]
  assign io_in_ready = _T_1390 | _T_1393; // @[IDU.scala 170:15]
  assign io_out_valid = io_in_valid; // @[IDU.scala 169:16]
  assign io_out_bits_cf_instr = io_in_bits_instr; // @[IDU.scala 171:18]
  assign io_out_bits_cf_pc = io_in_bits_pc; // @[IDU.scala 171:18]
  assign io_out_bits_cf_pnpc = io_in_bits_pnpc; // @[IDU.scala 171:18]
  assign io_out_bits_cf_exceptionVec_1 = _T_1423 & _T_1424; // @[IDU.scala 171:18 IDU.scala 185:37 IDU.scala 189:51]
  assign io_out_bits_cf_exceptionVec_2 = _T_1420 & io_in_valid; // @[IDU.scala 171:18 IDU.scala 185:37 IDU.scala 186:45]
  assign io_out_bits_cf_exceptionVec_12 = io_in_bits_exceptionVec_12; // @[IDU.scala 171:18 IDU.scala 185:37 IDU.scala 187:47]
  assign io_out_bits_cf_intrVec_0 = intrVecIDU[0]; // @[IDU.scala 171:18 IDU.scala 179:68]
  assign io_out_bits_cf_intrVec_1 = intrVecIDU[1]; // @[IDU.scala 171:18 IDU.scala 179:68]
  assign io_out_bits_cf_intrVec_2 = intrVecIDU[2]; // @[IDU.scala 171:18 IDU.scala 179:68]
  assign io_out_bits_cf_intrVec_3 = intrVecIDU[3]; // @[IDU.scala 171:18 IDU.scala 179:68]
  assign io_out_bits_cf_intrVec_4 = intrVecIDU[4]; // @[IDU.scala 171:18 IDU.scala 179:68]
  assign io_out_bits_cf_intrVec_5 = intrVecIDU[5]; // @[IDU.scala 171:18 IDU.scala 179:68]
  assign io_out_bits_cf_intrVec_6 = intrVecIDU[6]; // @[IDU.scala 171:18 IDU.scala 179:68]
  assign io_out_bits_cf_intrVec_7 = intrVecIDU[7]; // @[IDU.scala 171:18 IDU.scala 179:68]
  assign io_out_bits_cf_intrVec_8 = intrVecIDU[8]; // @[IDU.scala 171:18 IDU.scala 179:68]
  assign io_out_bits_cf_intrVec_9 = intrVecIDU[9]; // @[IDU.scala 171:18 IDU.scala 179:68]
  assign io_out_bits_cf_intrVec_10 = intrVecIDU[10]; // @[IDU.scala 171:18 IDU.scala 179:68]
  assign io_out_bits_cf_intrVec_11 = intrVecIDU[11]; // @[IDU.scala 171:18 IDU.scala 179:68]
  assign io_out_bits_cf_brIdx = io_in_bits_brIdx; // @[IDU.scala 171:18]
  assign io_out_bits_cf_crossPageIPFFix = io_in_bits_crossPageIPFFix; // @[IDU.scala 171:18]
  assign io_out_bits_ctrl_src1Type = {{1'd0}, _T_1379}; // @[IDU.scala 149:29]
  assign io_out_bits_ctrl_src2Type = {{1'd0}, src2Type}; // @[IDU.scala 150:29]
  assign io_out_bits_ctrl_fuType = _T_678 ? 3'h3 : decodeList_1; // @[IDU.scala 44:27]
  assign io_out_bits_ctrl_fuOpType = _T_1364 ? _GEN_3 : fuOpType; // @[IDU.scala 45:29 IDU.scala 142:85 IDU.scala 144:57 IDU.scala 145:57]
  assign io_out_bits_ctrl_rfSrc1 = src1Type ? 5'h0 : rfSrc1; // @[IDU.scala 97:27]
  assign io_out_bits_ctrl_rfSrc2 = _T_1087 ? rfSrc2 : 5'h0; // @[IDU.scala 98:27]
  assign io_out_bits_ctrl_rfWen = instrType[2]; // @[IDU.scala 99:27]
  assign io_out_bits_ctrl_rfDest = instrType[2] ? rfDest : 5'h0; // @[IDU.scala 100:27]
  assign io_out_bits_ctrl_isNutCoreTrap = _T_99 & io_in_valid; // @[IDU.scala 160:34 IDU.scala 194:34]
  assign io_out_bits_data_imm = isRVC ? immrvc : imm; // @[IDU.scala 138:25]
  assign io_isWFI = _T_203 & io_in_valid; // @[IDU.scala 195:12]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  _T_1396 = _RAND_0[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_1396 <= 64'h0;
    end else begin
      _T_1396 <= _T_1398;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1400 & _T_1402) begin
          $fwrite(32'h80000002,"[%d] Decoder: ",_T_1396); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1400 & _T_1402) begin
          $fwrite(32'h80000002,"issue: pc %x npc %x instr %x\n",io_out_bits_cf_pc,io_out_bits_cf_pnpc,io_out_bits_cf_instr); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Decoder_1(
  input         clock,
  input         reset,
  output        io_out_valid,
  output [63:0] io_out_bits_cf_instr,
  output [38:0] io_out_bits_cf_pc,
  output [38:0] io_out_bits_cf_pnpc,
  output        io_out_bits_cf_intrVec_0,
  output        io_out_bits_cf_intrVec_1,
  output        io_out_bits_cf_intrVec_2,
  output        io_out_bits_cf_intrVec_3,
  output        io_out_bits_cf_intrVec_4,
  output        io_out_bits_cf_intrVec_5,
  output        io_out_bits_cf_intrVec_6,
  output        io_out_bits_cf_intrVec_7,
  output        io_out_bits_cf_intrVec_8,
  output        io_out_bits_cf_intrVec_9,
  output        io_out_bits_cf_intrVec_10,
  output        io_out_bits_cf_intrVec_11,
  input         DISPLAY_ENABLE,
  input  [11:0] intrVecIDU
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] _T_1396; // @[GTimer.scala 24:20]
  wire [63:0] _T_1398 = _T_1396 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_1400 = io_out_valid & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  wire  _T_1402 = ~reset; // @[Debug.scala 56:24]
  assign io_out_valid = 1'h0; // @[IDU.scala 169:16]
  assign io_out_bits_cf_instr = 64'h0; // @[IDU.scala 171:18]
  assign io_out_bits_cf_pc = 39'h0; // @[IDU.scala 171:18]
  assign io_out_bits_cf_pnpc = 39'h0; // @[IDU.scala 171:18]
  assign io_out_bits_cf_intrVec_0 = intrVecIDU[0]; // @[IDU.scala 171:18 IDU.scala 179:68]
  assign io_out_bits_cf_intrVec_1 = intrVecIDU[1]; // @[IDU.scala 171:18 IDU.scala 179:68]
  assign io_out_bits_cf_intrVec_2 = intrVecIDU[2]; // @[IDU.scala 171:18 IDU.scala 179:68]
  assign io_out_bits_cf_intrVec_3 = intrVecIDU[3]; // @[IDU.scala 171:18 IDU.scala 179:68]
  assign io_out_bits_cf_intrVec_4 = intrVecIDU[4]; // @[IDU.scala 171:18 IDU.scala 179:68]
  assign io_out_bits_cf_intrVec_5 = intrVecIDU[5]; // @[IDU.scala 171:18 IDU.scala 179:68]
  assign io_out_bits_cf_intrVec_6 = intrVecIDU[6]; // @[IDU.scala 171:18 IDU.scala 179:68]
  assign io_out_bits_cf_intrVec_7 = intrVecIDU[7]; // @[IDU.scala 171:18 IDU.scala 179:68]
  assign io_out_bits_cf_intrVec_8 = intrVecIDU[8]; // @[IDU.scala 171:18 IDU.scala 179:68]
  assign io_out_bits_cf_intrVec_9 = intrVecIDU[9]; // @[IDU.scala 171:18 IDU.scala 179:68]
  assign io_out_bits_cf_intrVec_10 = intrVecIDU[10]; // @[IDU.scala 171:18 IDU.scala 179:68]
  assign io_out_bits_cf_intrVec_11 = intrVecIDU[11]; // @[IDU.scala 171:18 IDU.scala 179:68]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  _T_1396 = _RAND_0[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_1396 <= 64'h0;
    end else begin
      _T_1396 <= _T_1398;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1400 & _T_1402) begin
          $fwrite(32'h80000002,"[%d] Decoder_1: ",_T_1396); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1400 & _T_1402) begin
          $fwrite(32'h80000002,"issue: pc %x npc %x instr %x\n",io_out_bits_cf_pc,io_out_bits_cf_pnpc,io_out_bits_cf_instr); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module IDU(
  input         clock,
  input         reset,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [63:0] io_in_0_bits_instr,
  input  [38:0] io_in_0_bits_pc,
  input  [38:0] io_in_0_bits_pnpc,
  input         io_in_0_bits_exceptionVec_12,
  input  [3:0]  io_in_0_bits_brIdx,
  input         io_in_0_bits_crossPageIPFFix,
  input         io_out_0_ready,
  output        io_out_0_valid,
  output [63:0] io_out_0_bits_cf_instr,
  output [38:0] io_out_0_bits_cf_pc,
  output [38:0] io_out_0_bits_cf_pnpc,
  output        io_out_0_bits_cf_exceptionVec_1,
  output        io_out_0_bits_cf_exceptionVec_2,
  output        io_out_0_bits_cf_exceptionVec_12,
  output        io_out_0_bits_cf_intrVec_0,
  output        io_out_0_bits_cf_intrVec_1,
  output        io_out_0_bits_cf_intrVec_2,
  output        io_out_0_bits_cf_intrVec_3,
  output        io_out_0_bits_cf_intrVec_4,
  output        io_out_0_bits_cf_intrVec_5,
  output        io_out_0_bits_cf_intrVec_6,
  output        io_out_0_bits_cf_intrVec_7,
  output        io_out_0_bits_cf_intrVec_8,
  output        io_out_0_bits_cf_intrVec_9,
  output        io_out_0_bits_cf_intrVec_10,
  output        io_out_0_bits_cf_intrVec_11,
  output [3:0]  io_out_0_bits_cf_brIdx,
  output        io_out_0_bits_cf_crossPageIPFFix,
  output [1:0]  io_out_0_bits_ctrl_src1Type,
  output [1:0]  io_out_0_bits_ctrl_src2Type,
  output [2:0]  io_out_0_bits_ctrl_fuType,
  output [6:0]  io_out_0_bits_ctrl_fuOpType,
  output [4:0]  io_out_0_bits_ctrl_rfSrc1,
  output [4:0]  io_out_0_bits_ctrl_rfSrc2,
  output        io_out_0_bits_ctrl_rfWen,
  output [4:0]  io_out_0_bits_ctrl_rfDest,
  output        io_out_0_bits_ctrl_isNutCoreTrap,
  output [63:0] io_out_0_bits_data_imm,
  output        io_out_1_bits_cf_intrVec_0,
  output        io_out_1_bits_cf_intrVec_1,
  output        io_out_1_bits_cf_intrVec_2,
  output        io_out_1_bits_cf_intrVec_3,
  output        io_out_1_bits_cf_intrVec_4,
  output        io_out_1_bits_cf_intrVec_5,
  output        io_out_1_bits_cf_intrVec_6,
  output        io_out_1_bits_cf_intrVec_7,
  output        io_out_1_bits_cf_intrVec_8,
  output        io_out_1_bits_cf_intrVec_9,
  output        io_out_1_bits_cf_intrVec_10,
  output        io_out_1_bits_cf_intrVec_11,
  input         _T_13,
  input         vmEnable,
  input  [11:0] intrVec,
  output        _T_0
);
  wire  decoder1_clock; // @[IDU.scala 204:25]
  wire  decoder1_reset; // @[IDU.scala 204:25]
  wire  decoder1_io_in_ready; // @[IDU.scala 204:25]
  wire  decoder1_io_in_valid; // @[IDU.scala 204:25]
  wire [63:0] decoder1_io_in_bits_instr; // @[IDU.scala 204:25]
  wire [38:0] decoder1_io_in_bits_pc; // @[IDU.scala 204:25]
  wire [38:0] decoder1_io_in_bits_pnpc; // @[IDU.scala 204:25]
  wire  decoder1_io_in_bits_exceptionVec_12; // @[IDU.scala 204:25]
  wire [3:0] decoder1_io_in_bits_brIdx; // @[IDU.scala 204:25]
  wire  decoder1_io_in_bits_crossPageIPFFix; // @[IDU.scala 204:25]
  wire  decoder1_io_out_ready; // @[IDU.scala 204:25]
  wire  decoder1_io_out_valid; // @[IDU.scala 204:25]
  wire [63:0] decoder1_io_out_bits_cf_instr; // @[IDU.scala 204:25]
  wire [38:0] decoder1_io_out_bits_cf_pc; // @[IDU.scala 204:25]
  wire [38:0] decoder1_io_out_bits_cf_pnpc; // @[IDU.scala 204:25]
  wire  decoder1_io_out_bits_cf_exceptionVec_1; // @[IDU.scala 204:25]
  wire  decoder1_io_out_bits_cf_exceptionVec_2; // @[IDU.scala 204:25]
  wire  decoder1_io_out_bits_cf_exceptionVec_12; // @[IDU.scala 204:25]
  wire  decoder1_io_out_bits_cf_intrVec_0; // @[IDU.scala 204:25]
  wire  decoder1_io_out_bits_cf_intrVec_1; // @[IDU.scala 204:25]
  wire  decoder1_io_out_bits_cf_intrVec_2; // @[IDU.scala 204:25]
  wire  decoder1_io_out_bits_cf_intrVec_3; // @[IDU.scala 204:25]
  wire  decoder1_io_out_bits_cf_intrVec_4; // @[IDU.scala 204:25]
  wire  decoder1_io_out_bits_cf_intrVec_5; // @[IDU.scala 204:25]
  wire  decoder1_io_out_bits_cf_intrVec_6; // @[IDU.scala 204:25]
  wire  decoder1_io_out_bits_cf_intrVec_7; // @[IDU.scala 204:25]
  wire  decoder1_io_out_bits_cf_intrVec_8; // @[IDU.scala 204:25]
  wire  decoder1_io_out_bits_cf_intrVec_9; // @[IDU.scala 204:25]
  wire  decoder1_io_out_bits_cf_intrVec_10; // @[IDU.scala 204:25]
  wire  decoder1_io_out_bits_cf_intrVec_11; // @[IDU.scala 204:25]
  wire [3:0] decoder1_io_out_bits_cf_brIdx; // @[IDU.scala 204:25]
  wire  decoder1_io_out_bits_cf_crossPageIPFFix; // @[IDU.scala 204:25]
  wire [1:0] decoder1_io_out_bits_ctrl_src1Type; // @[IDU.scala 204:25]
  wire [1:0] decoder1_io_out_bits_ctrl_src2Type; // @[IDU.scala 204:25]
  wire [2:0] decoder1_io_out_bits_ctrl_fuType; // @[IDU.scala 204:25]
  wire [6:0] decoder1_io_out_bits_ctrl_fuOpType; // @[IDU.scala 204:25]
  wire [4:0] decoder1_io_out_bits_ctrl_rfSrc1; // @[IDU.scala 204:25]
  wire [4:0] decoder1_io_out_bits_ctrl_rfSrc2; // @[IDU.scala 204:25]
  wire  decoder1_io_out_bits_ctrl_rfWen; // @[IDU.scala 204:25]
  wire [4:0] decoder1_io_out_bits_ctrl_rfDest; // @[IDU.scala 204:25]
  wire  decoder1_io_out_bits_ctrl_isNutCoreTrap; // @[IDU.scala 204:25]
  wire [63:0] decoder1_io_out_bits_data_imm; // @[IDU.scala 204:25]
  wire  decoder1_io_isWFI; // @[IDU.scala 204:25]
  wire  decoder1_DISPLAY_ENABLE; // @[IDU.scala 204:25]
  wire  decoder1_DTLBENABLE; // @[IDU.scala 204:25]
  wire [11:0] decoder1_intrVecIDU; // @[IDU.scala 204:25]
  wire  decoder2_clock; // @[IDU.scala 205:25]
  wire  decoder2_reset; // @[IDU.scala 205:25]
  wire  decoder2_io_out_valid; // @[IDU.scala 205:25]
  wire [63:0] decoder2_io_out_bits_cf_instr; // @[IDU.scala 205:25]
  wire [38:0] decoder2_io_out_bits_cf_pc; // @[IDU.scala 205:25]
  wire [38:0] decoder2_io_out_bits_cf_pnpc; // @[IDU.scala 205:25]
  wire  decoder2_io_out_bits_cf_intrVec_0; // @[IDU.scala 205:25]
  wire  decoder2_io_out_bits_cf_intrVec_1; // @[IDU.scala 205:25]
  wire  decoder2_io_out_bits_cf_intrVec_2; // @[IDU.scala 205:25]
  wire  decoder2_io_out_bits_cf_intrVec_3; // @[IDU.scala 205:25]
  wire  decoder2_io_out_bits_cf_intrVec_4; // @[IDU.scala 205:25]
  wire  decoder2_io_out_bits_cf_intrVec_5; // @[IDU.scala 205:25]
  wire  decoder2_io_out_bits_cf_intrVec_6; // @[IDU.scala 205:25]
  wire  decoder2_io_out_bits_cf_intrVec_7; // @[IDU.scala 205:25]
  wire  decoder2_io_out_bits_cf_intrVec_8; // @[IDU.scala 205:25]
  wire  decoder2_io_out_bits_cf_intrVec_9; // @[IDU.scala 205:25]
  wire  decoder2_io_out_bits_cf_intrVec_10; // @[IDU.scala 205:25]
  wire  decoder2_io_out_bits_cf_intrVec_11; // @[IDU.scala 205:25]
  wire  decoder2_DISPLAY_ENABLE; // @[IDU.scala 205:25]
  wire [11:0] decoder2_intrVecIDU; // @[IDU.scala 205:25]
  wire  _T = decoder1_io_isWFI; // @[IDU.scala 216:45]
  Decoder decoder1 ( // @[IDU.scala 204:25]
    .clock(decoder1_clock),
    .reset(decoder1_reset),
    .io_in_ready(decoder1_io_in_ready),
    .io_in_valid(decoder1_io_in_valid),
    .io_in_bits_instr(decoder1_io_in_bits_instr),
    .io_in_bits_pc(decoder1_io_in_bits_pc),
    .io_in_bits_pnpc(decoder1_io_in_bits_pnpc),
    .io_in_bits_exceptionVec_12(decoder1_io_in_bits_exceptionVec_12),
    .io_in_bits_brIdx(decoder1_io_in_bits_brIdx),
    .io_in_bits_crossPageIPFFix(decoder1_io_in_bits_crossPageIPFFix),
    .io_out_ready(decoder1_io_out_ready),
    .io_out_valid(decoder1_io_out_valid),
    .io_out_bits_cf_instr(decoder1_io_out_bits_cf_instr),
    .io_out_bits_cf_pc(decoder1_io_out_bits_cf_pc),
    .io_out_bits_cf_pnpc(decoder1_io_out_bits_cf_pnpc),
    .io_out_bits_cf_exceptionVec_1(decoder1_io_out_bits_cf_exceptionVec_1),
    .io_out_bits_cf_exceptionVec_2(decoder1_io_out_bits_cf_exceptionVec_2),
    .io_out_bits_cf_exceptionVec_12(decoder1_io_out_bits_cf_exceptionVec_12),
    .io_out_bits_cf_intrVec_0(decoder1_io_out_bits_cf_intrVec_0),
    .io_out_bits_cf_intrVec_1(decoder1_io_out_bits_cf_intrVec_1),
    .io_out_bits_cf_intrVec_2(decoder1_io_out_bits_cf_intrVec_2),
    .io_out_bits_cf_intrVec_3(decoder1_io_out_bits_cf_intrVec_3),
    .io_out_bits_cf_intrVec_4(decoder1_io_out_bits_cf_intrVec_4),
    .io_out_bits_cf_intrVec_5(decoder1_io_out_bits_cf_intrVec_5),
    .io_out_bits_cf_intrVec_6(decoder1_io_out_bits_cf_intrVec_6),
    .io_out_bits_cf_intrVec_7(decoder1_io_out_bits_cf_intrVec_7),
    .io_out_bits_cf_intrVec_8(decoder1_io_out_bits_cf_intrVec_8),
    .io_out_bits_cf_intrVec_9(decoder1_io_out_bits_cf_intrVec_9),
    .io_out_bits_cf_intrVec_10(decoder1_io_out_bits_cf_intrVec_10),
    .io_out_bits_cf_intrVec_11(decoder1_io_out_bits_cf_intrVec_11),
    .io_out_bits_cf_brIdx(decoder1_io_out_bits_cf_brIdx),
    .io_out_bits_cf_crossPageIPFFix(decoder1_io_out_bits_cf_crossPageIPFFix),
    .io_out_bits_ctrl_src1Type(decoder1_io_out_bits_ctrl_src1Type),
    .io_out_bits_ctrl_src2Type(decoder1_io_out_bits_ctrl_src2Type),
    .io_out_bits_ctrl_fuType(decoder1_io_out_bits_ctrl_fuType),
    .io_out_bits_ctrl_fuOpType(decoder1_io_out_bits_ctrl_fuOpType),
    .io_out_bits_ctrl_rfSrc1(decoder1_io_out_bits_ctrl_rfSrc1),
    .io_out_bits_ctrl_rfSrc2(decoder1_io_out_bits_ctrl_rfSrc2),
    .io_out_bits_ctrl_rfWen(decoder1_io_out_bits_ctrl_rfWen),
    .io_out_bits_ctrl_rfDest(decoder1_io_out_bits_ctrl_rfDest),
    .io_out_bits_ctrl_isNutCoreTrap(decoder1_io_out_bits_ctrl_isNutCoreTrap),
    .io_out_bits_data_imm(decoder1_io_out_bits_data_imm),
    .io_isWFI(decoder1_io_isWFI),
    .DISPLAY_ENABLE(decoder1_DISPLAY_ENABLE),
    .DTLBENABLE(decoder1_DTLBENABLE),
    .intrVecIDU(decoder1_intrVecIDU)
  );
  Decoder_1 decoder2 ( // @[IDU.scala 205:25]
    .clock(decoder2_clock),
    .reset(decoder2_reset),
    .io_out_valid(decoder2_io_out_valid),
    .io_out_bits_cf_instr(decoder2_io_out_bits_cf_instr),
    .io_out_bits_cf_pc(decoder2_io_out_bits_cf_pc),
    .io_out_bits_cf_pnpc(decoder2_io_out_bits_cf_pnpc),
    .io_out_bits_cf_intrVec_0(decoder2_io_out_bits_cf_intrVec_0),
    .io_out_bits_cf_intrVec_1(decoder2_io_out_bits_cf_intrVec_1),
    .io_out_bits_cf_intrVec_2(decoder2_io_out_bits_cf_intrVec_2),
    .io_out_bits_cf_intrVec_3(decoder2_io_out_bits_cf_intrVec_3),
    .io_out_bits_cf_intrVec_4(decoder2_io_out_bits_cf_intrVec_4),
    .io_out_bits_cf_intrVec_5(decoder2_io_out_bits_cf_intrVec_5),
    .io_out_bits_cf_intrVec_6(decoder2_io_out_bits_cf_intrVec_6),
    .io_out_bits_cf_intrVec_7(decoder2_io_out_bits_cf_intrVec_7),
    .io_out_bits_cf_intrVec_8(decoder2_io_out_bits_cf_intrVec_8),
    .io_out_bits_cf_intrVec_9(decoder2_io_out_bits_cf_intrVec_9),
    .io_out_bits_cf_intrVec_10(decoder2_io_out_bits_cf_intrVec_10),
    .io_out_bits_cf_intrVec_11(decoder2_io_out_bits_cf_intrVec_11),
    .DISPLAY_ENABLE(decoder2_DISPLAY_ENABLE),
    .intrVecIDU(decoder2_intrVecIDU)
  );
  assign io_in_0_ready = decoder1_io_in_ready; // @[IDU.scala 206:12]
  assign io_out_0_valid = decoder1_io_out_valid; // @[IDU.scala 208:13]
  assign io_out_0_bits_cf_instr = decoder1_io_out_bits_cf_instr; // @[IDU.scala 208:13]
  assign io_out_0_bits_cf_pc = decoder1_io_out_bits_cf_pc; // @[IDU.scala 208:13]
  assign io_out_0_bits_cf_pnpc = decoder1_io_out_bits_cf_pnpc; // @[IDU.scala 208:13]
  assign io_out_0_bits_cf_exceptionVec_1 = decoder1_io_out_bits_cf_exceptionVec_1; // @[IDU.scala 208:13]
  assign io_out_0_bits_cf_exceptionVec_2 = decoder1_io_out_bits_cf_exceptionVec_2; // @[IDU.scala 208:13]
  assign io_out_0_bits_cf_exceptionVec_12 = decoder1_io_out_bits_cf_exceptionVec_12; // @[IDU.scala 208:13]
  assign io_out_0_bits_cf_intrVec_0 = decoder1_io_out_bits_cf_intrVec_0; // @[IDU.scala 208:13]
  assign io_out_0_bits_cf_intrVec_1 = decoder1_io_out_bits_cf_intrVec_1; // @[IDU.scala 208:13]
  assign io_out_0_bits_cf_intrVec_2 = decoder1_io_out_bits_cf_intrVec_2; // @[IDU.scala 208:13]
  assign io_out_0_bits_cf_intrVec_3 = decoder1_io_out_bits_cf_intrVec_3; // @[IDU.scala 208:13]
  assign io_out_0_bits_cf_intrVec_4 = decoder1_io_out_bits_cf_intrVec_4; // @[IDU.scala 208:13]
  assign io_out_0_bits_cf_intrVec_5 = decoder1_io_out_bits_cf_intrVec_5; // @[IDU.scala 208:13]
  assign io_out_0_bits_cf_intrVec_6 = decoder1_io_out_bits_cf_intrVec_6; // @[IDU.scala 208:13]
  assign io_out_0_bits_cf_intrVec_7 = decoder1_io_out_bits_cf_intrVec_7; // @[IDU.scala 208:13]
  assign io_out_0_bits_cf_intrVec_8 = decoder1_io_out_bits_cf_intrVec_8; // @[IDU.scala 208:13]
  assign io_out_0_bits_cf_intrVec_9 = decoder1_io_out_bits_cf_intrVec_9; // @[IDU.scala 208:13]
  assign io_out_0_bits_cf_intrVec_10 = decoder1_io_out_bits_cf_intrVec_10; // @[IDU.scala 208:13]
  assign io_out_0_bits_cf_intrVec_11 = decoder1_io_out_bits_cf_intrVec_11; // @[IDU.scala 208:13]
  assign io_out_0_bits_cf_brIdx = decoder1_io_out_bits_cf_brIdx; // @[IDU.scala 208:13]
  assign io_out_0_bits_cf_crossPageIPFFix = decoder1_io_out_bits_cf_crossPageIPFFix; // @[IDU.scala 208:13]
  assign io_out_0_bits_ctrl_src1Type = decoder1_io_out_bits_ctrl_src1Type; // @[IDU.scala 208:13]
  assign io_out_0_bits_ctrl_src2Type = decoder1_io_out_bits_ctrl_src2Type; // @[IDU.scala 208:13]
  assign io_out_0_bits_ctrl_fuType = decoder1_io_out_bits_ctrl_fuType; // @[IDU.scala 208:13]
  assign io_out_0_bits_ctrl_fuOpType = decoder1_io_out_bits_ctrl_fuOpType; // @[IDU.scala 208:13]
  assign io_out_0_bits_ctrl_rfSrc1 = decoder1_io_out_bits_ctrl_rfSrc1; // @[IDU.scala 208:13]
  assign io_out_0_bits_ctrl_rfSrc2 = decoder1_io_out_bits_ctrl_rfSrc2; // @[IDU.scala 208:13]
  assign io_out_0_bits_ctrl_rfWen = decoder1_io_out_bits_ctrl_rfWen; // @[IDU.scala 208:13]
  assign io_out_0_bits_ctrl_rfDest = decoder1_io_out_bits_ctrl_rfDest; // @[IDU.scala 208:13]
  assign io_out_0_bits_ctrl_isNutCoreTrap = decoder1_io_out_bits_ctrl_isNutCoreTrap; // @[IDU.scala 208:13]
  assign io_out_0_bits_data_imm = decoder1_io_out_bits_data_imm; // @[IDU.scala 208:13]
  assign io_out_1_bits_cf_intrVec_0 = decoder2_io_out_bits_cf_intrVec_0; // @[IDU.scala 209:13]
  assign io_out_1_bits_cf_intrVec_1 = decoder2_io_out_bits_cf_intrVec_1; // @[IDU.scala 209:13]
  assign io_out_1_bits_cf_intrVec_2 = decoder2_io_out_bits_cf_intrVec_2; // @[IDU.scala 209:13]
  assign io_out_1_bits_cf_intrVec_3 = decoder2_io_out_bits_cf_intrVec_3; // @[IDU.scala 209:13]
  assign io_out_1_bits_cf_intrVec_4 = decoder2_io_out_bits_cf_intrVec_4; // @[IDU.scala 209:13]
  assign io_out_1_bits_cf_intrVec_5 = decoder2_io_out_bits_cf_intrVec_5; // @[IDU.scala 209:13]
  assign io_out_1_bits_cf_intrVec_6 = decoder2_io_out_bits_cf_intrVec_6; // @[IDU.scala 209:13]
  assign io_out_1_bits_cf_intrVec_7 = decoder2_io_out_bits_cf_intrVec_7; // @[IDU.scala 209:13]
  assign io_out_1_bits_cf_intrVec_8 = decoder2_io_out_bits_cf_intrVec_8; // @[IDU.scala 209:13]
  assign io_out_1_bits_cf_intrVec_9 = decoder2_io_out_bits_cf_intrVec_9; // @[IDU.scala 209:13]
  assign io_out_1_bits_cf_intrVec_10 = decoder2_io_out_bits_cf_intrVec_10; // @[IDU.scala 209:13]
  assign io_out_1_bits_cf_intrVec_11 = decoder2_io_out_bits_cf_intrVec_11; // @[IDU.scala 209:13]
  assign _T_0 = _T;
  assign decoder1_clock = clock;
  assign decoder1_reset = reset;
  assign decoder1_io_in_valid = io_in_0_valid; // @[IDU.scala 206:12]
  assign decoder1_io_in_bits_instr = io_in_0_bits_instr; // @[IDU.scala 206:12]
  assign decoder1_io_in_bits_pc = io_in_0_bits_pc; // @[IDU.scala 206:12]
  assign decoder1_io_in_bits_pnpc = io_in_0_bits_pnpc; // @[IDU.scala 206:12]
  assign decoder1_io_in_bits_exceptionVec_12 = io_in_0_bits_exceptionVec_12; // @[IDU.scala 206:12]
  assign decoder1_io_in_bits_brIdx = io_in_0_bits_brIdx; // @[IDU.scala 206:12]
  assign decoder1_io_in_bits_crossPageIPFFix = io_in_0_bits_crossPageIPFFix; // @[IDU.scala 206:12]
  assign decoder1_io_out_ready = io_out_0_ready; // @[IDU.scala 208:13]
  assign decoder1_DISPLAY_ENABLE = _T_13;
  assign decoder1_DTLBENABLE = vmEnable;
  assign decoder1_intrVecIDU = intrVec;
  assign decoder2_clock = clock;
  assign decoder2_reset = reset;
  assign decoder2_DISPLAY_ENABLE = _T_13;
  assign decoder2_intrVecIDU = intrVec;
endmodule
module FlushableQueue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits_instr,
  input  [38:0] io_enq_bits_pc,
  input  [38:0] io_enq_bits_pnpc,
  input         io_enq_bits_exceptionVec_12,
  input  [3:0]  io_enq_bits_brIdx,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits_instr,
  output [38:0] io_deq_bits_pc,
  output [38:0] io_deq_bits_pnpc,
  output        io_deq_bits_exceptionVec_12,
  output [3:0]  io_deq_bits_brIdx,
  input         io_flush
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram_instr [0:3]; // @[FlushableQueue.scala 33:24]
  wire [63:0] ram_instr__T_15_data; // @[FlushableQueue.scala 33:24]
  wire [1:0] ram_instr__T_15_addr; // @[FlushableQueue.scala 33:24]
  wire [63:0] ram_instr__T_5_data; // @[FlushableQueue.scala 33:24]
  wire [1:0] ram_instr__T_5_addr; // @[FlushableQueue.scala 33:24]
  wire  ram_instr__T_5_mask; // @[FlushableQueue.scala 33:24]
  wire  ram_instr__T_5_en; // @[FlushableQueue.scala 33:24]
  reg [38:0] ram_pc [0:3]; // @[FlushableQueue.scala 33:24]
  wire [38:0] ram_pc__T_15_data; // @[FlushableQueue.scala 33:24]
  wire [1:0] ram_pc__T_15_addr; // @[FlushableQueue.scala 33:24]
  wire [38:0] ram_pc__T_5_data; // @[FlushableQueue.scala 33:24]
  wire [1:0] ram_pc__T_5_addr; // @[FlushableQueue.scala 33:24]
  wire  ram_pc__T_5_mask; // @[FlushableQueue.scala 33:24]
  wire  ram_pc__T_5_en; // @[FlushableQueue.scala 33:24]
  reg [38:0] ram_pnpc [0:3]; // @[FlushableQueue.scala 33:24]
  wire [38:0] ram_pnpc__T_15_data; // @[FlushableQueue.scala 33:24]
  wire [1:0] ram_pnpc__T_15_addr; // @[FlushableQueue.scala 33:24]
  wire [38:0] ram_pnpc__T_5_data; // @[FlushableQueue.scala 33:24]
  wire [1:0] ram_pnpc__T_5_addr; // @[FlushableQueue.scala 33:24]
  wire  ram_pnpc__T_5_mask; // @[FlushableQueue.scala 33:24]
  wire  ram_pnpc__T_5_en; // @[FlushableQueue.scala 33:24]
  reg  ram_exceptionVec_12 [0:3]; // @[FlushableQueue.scala 33:24]
  wire  ram_exceptionVec_12__T_15_data; // @[FlushableQueue.scala 33:24]
  wire [1:0] ram_exceptionVec_12__T_15_addr; // @[FlushableQueue.scala 33:24]
  wire  ram_exceptionVec_12__T_5_data; // @[FlushableQueue.scala 33:24]
  wire [1:0] ram_exceptionVec_12__T_5_addr; // @[FlushableQueue.scala 33:24]
  wire  ram_exceptionVec_12__T_5_mask; // @[FlushableQueue.scala 33:24]
  wire  ram_exceptionVec_12__T_5_en; // @[FlushableQueue.scala 33:24]
  reg [3:0] ram_brIdx [0:3]; // @[FlushableQueue.scala 33:24]
  wire [3:0] ram_brIdx__T_15_data; // @[FlushableQueue.scala 33:24]
  wire [1:0] ram_brIdx__T_15_addr; // @[FlushableQueue.scala 33:24]
  wire [3:0] ram_brIdx__T_5_data; // @[FlushableQueue.scala 33:24]
  wire [1:0] ram_brIdx__T_5_addr; // @[FlushableQueue.scala 33:24]
  wire  ram_brIdx__T_5_mask; // @[FlushableQueue.scala 33:24]
  wire  ram_brIdx__T_5_en; // @[FlushableQueue.scala 33:24]
  reg [1:0] value; // @[Counter.scala 29:33]
  reg [1:0] value_1; // @[Counter.scala 29:33]
  reg  maybe_full; // @[FlushableQueue.scala 36:35]
  wire  _T = value == value_1; // @[FlushableQueue.scala 38:41]
  wire  _T_1 = ~maybe_full; // @[FlushableQueue.scala 39:36]
  wire  empty = _T & _T_1; // @[FlushableQueue.scala 39:33]
  wire  _T_2 = _T & maybe_full; // @[FlushableQueue.scala 40:32]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _T_8 = value + 2'h1; // @[Counter.scala 39:22]
  wire [1:0] _T_11 = value_1 + 2'h1; // @[Counter.scala 39:22]
  wire  _T_12 = do_enq != do_deq; // @[FlushableQueue.scala 51:16]
  assign ram_instr__T_15_addr = value_1;
  assign ram_instr__T_15_data = ram_instr[ram_instr__T_15_addr]; // @[FlushableQueue.scala 33:24]
  assign ram_instr__T_5_data = io_enq_bits_instr;
  assign ram_instr__T_5_addr = value;
  assign ram_instr__T_5_mask = 1'h1;
  assign ram_instr__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_pc__T_15_addr = value_1;
  assign ram_pc__T_15_data = ram_pc[ram_pc__T_15_addr]; // @[FlushableQueue.scala 33:24]
  assign ram_pc__T_5_data = io_enq_bits_pc;
  assign ram_pc__T_5_addr = value;
  assign ram_pc__T_5_mask = 1'h1;
  assign ram_pc__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_pnpc__T_15_addr = value_1;
  assign ram_pnpc__T_15_data = ram_pnpc[ram_pnpc__T_15_addr]; // @[FlushableQueue.scala 33:24]
  assign ram_pnpc__T_5_data = io_enq_bits_pnpc;
  assign ram_pnpc__T_5_addr = value;
  assign ram_pnpc__T_5_mask = 1'h1;
  assign ram_pnpc__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_12__T_15_addr = value_1;
  assign ram_exceptionVec_12__T_15_data = ram_exceptionVec_12[ram_exceptionVec_12__T_15_addr]; // @[FlushableQueue.scala 33:24]
  assign ram_exceptionVec_12__T_5_data = io_enq_bits_exceptionVec_12;
  assign ram_exceptionVec_12__T_5_addr = value;
  assign ram_exceptionVec_12__T_5_mask = 1'h1;
  assign ram_exceptionVec_12__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_brIdx__T_15_addr = value_1;
  assign ram_brIdx__T_15_data = ram_brIdx[ram_brIdx__T_15_addr]; // @[FlushableQueue.scala 33:24]
  assign ram_brIdx__T_5_data = io_enq_bits_brIdx;
  assign ram_brIdx__T_5_addr = value;
  assign ram_brIdx__T_5_mask = 1'h1;
  assign ram_brIdx__T_5_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~_T_2; // @[FlushableQueue.scala 56:16]
  assign io_deq_valid = ~empty; // @[FlushableQueue.scala 55:16]
  assign io_deq_bits_instr = ram_instr__T_15_data; // @[FlushableQueue.scala 57:15]
  assign io_deq_bits_pc = ram_pc__T_15_data; // @[FlushableQueue.scala 57:15]
  assign io_deq_bits_pnpc = ram_pnpc__T_15_data; // @[FlushableQueue.scala 57:15]
  assign io_deq_bits_exceptionVec_12 = ram_exceptionVec_12__T_15_data; // @[FlushableQueue.scala 57:15]
  assign io_deq_bits_brIdx = ram_brIdx__T_15_data; // @[FlushableQueue.scala 57:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_instr[initvar] = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_pc[initvar] = _RAND_1[38:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_pnpc[initvar] = _RAND_2[38:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_12[initvar] = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_brIdx[initvar] = _RAND_4[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  value_1 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  maybe_full = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram_instr__T_5_en & ram_instr__T_5_mask) begin
      ram_instr[ram_instr__T_5_addr] <= ram_instr__T_5_data; // @[FlushableQueue.scala 33:24]
    end
    if(ram_pc__T_5_en & ram_pc__T_5_mask) begin
      ram_pc[ram_pc__T_5_addr] <= ram_pc__T_5_data; // @[FlushableQueue.scala 33:24]
    end
    if(ram_pnpc__T_5_en & ram_pnpc__T_5_mask) begin
      ram_pnpc[ram_pnpc__T_5_addr] <= ram_pnpc__T_5_data; // @[FlushableQueue.scala 33:24]
    end
    if(ram_exceptionVec_12__T_5_en & ram_exceptionVec_12__T_5_mask) begin
      ram_exceptionVec_12[ram_exceptionVec_12__T_5_addr] <= ram_exceptionVec_12__T_5_data; // @[FlushableQueue.scala 33:24]
    end
    if(ram_brIdx__T_5_en & ram_brIdx__T_5_mask) begin
      ram_brIdx[ram_brIdx__T_5_addr] <= ram_brIdx__T_5_data; // @[FlushableQueue.scala 33:24]
    end
    if (reset) begin
      value <= 2'h0;
    end else if (io_flush) begin
      value <= 2'h0;
    end else if (do_enq) begin
      value <= _T_8;
    end
    if (reset) begin
      value_1 <= 2'h0;
    end else if (io_flush) begin
      value_1 <= 2'h0;
    end else if (do_deq) begin
      value_1 <= _T_11;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else if (io_flush) begin
      maybe_full <= 1'h0;
    end else if (_T_12) begin
      maybe_full <= do_enq;
    end
  end
endmodule
module Frontend_inorder(
  input         clock,
  input         reset,
  input         io_out_0_ready,
  output        io_out_0_valid,
  output [63:0] io_out_0_bits_cf_instr,
  output [38:0] io_out_0_bits_cf_pc,
  output [38:0] io_out_0_bits_cf_pnpc,
  output        io_out_0_bits_cf_exceptionVec_1,
  output        io_out_0_bits_cf_exceptionVec_2,
  output        io_out_0_bits_cf_exceptionVec_12,
  output        io_out_0_bits_cf_intrVec_0,
  output        io_out_0_bits_cf_intrVec_1,
  output        io_out_0_bits_cf_intrVec_2,
  output        io_out_0_bits_cf_intrVec_3,
  output        io_out_0_bits_cf_intrVec_4,
  output        io_out_0_bits_cf_intrVec_5,
  output        io_out_0_bits_cf_intrVec_6,
  output        io_out_0_bits_cf_intrVec_7,
  output        io_out_0_bits_cf_intrVec_8,
  output        io_out_0_bits_cf_intrVec_9,
  output        io_out_0_bits_cf_intrVec_10,
  output        io_out_0_bits_cf_intrVec_11,
  output [3:0]  io_out_0_bits_cf_brIdx,
  output        io_out_0_bits_cf_crossPageIPFFix,
  output [1:0]  io_out_0_bits_ctrl_src1Type,
  output [1:0]  io_out_0_bits_ctrl_src2Type,
  output [2:0]  io_out_0_bits_ctrl_fuType,
  output [6:0]  io_out_0_bits_ctrl_fuOpType,
  output [4:0]  io_out_0_bits_ctrl_rfSrc1,
  output [4:0]  io_out_0_bits_ctrl_rfSrc2,
  output        io_out_0_bits_ctrl_rfWen,
  output [4:0]  io_out_0_bits_ctrl_rfDest,
  output        io_out_0_bits_ctrl_isNutCoreTrap,
  output [63:0] io_out_0_bits_data_imm,
  output        io_out_1_bits_cf_intrVec_0,
  output        io_out_1_bits_cf_intrVec_1,
  output        io_out_1_bits_cf_intrVec_2,
  output        io_out_1_bits_cf_intrVec_3,
  output        io_out_1_bits_cf_intrVec_4,
  output        io_out_1_bits_cf_intrVec_5,
  output        io_out_1_bits_cf_intrVec_6,
  output        io_out_1_bits_cf_intrVec_7,
  output        io_out_1_bits_cf_intrVec_8,
  output        io_out_1_bits_cf_intrVec_9,
  output        io_out_1_bits_cf_intrVec_10,
  output        io_out_1_bits_cf_intrVec_11,
  input         io_imem_req_ready,
  output        io_imem_req_valid,
  output [38:0] io_imem_req_bits_addr,
  output [86:0] io_imem_req_bits_user,
  output        io_imem_resp_ready,
  input         io_imem_resp_valid,
  input  [63:0] io_imem_resp_bits_rdata,
  input  [86:0] io_imem_resp_bits_user,
  output [3:0]  io_flushVec,
  input         io_ipf,
  input  [38:0] io_redirect_target,
  input         io_redirect_valid,
  input         flushICache,
  input         _T_243_valid,
  input  [38:0] _T_243_pc,
  input         _T_243_isMissPredict,
  input  [38:0] _T_243_actualTarget,
  input         _T_243_actualTaken,
  input  [6:0]  _T_243_fuOpType,
  input  [1:0]  _T_243_btbType,
  input         _T_243_isRVC,
  input         DISPLAY_ENABLE,
  input         vmEnable,
  input  [11:0] intrVec,
  output        _T_0,
  output        _T_65,
  input         flushTLB,
  output        _T_66
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire  ifu_clock; // @[Frontend.scala 106:20]
  wire  ifu_reset; // @[Frontend.scala 106:20]
  wire  ifu_io_imem_req_ready; // @[Frontend.scala 106:20]
  wire  ifu_io_imem_req_valid; // @[Frontend.scala 106:20]
  wire [38:0] ifu_io_imem_req_bits_addr; // @[Frontend.scala 106:20]
  wire [81:0] ifu_io_imem_req_bits_user; // @[Frontend.scala 106:20]
  wire  ifu_io_imem_resp_ready; // @[Frontend.scala 106:20]
  wire  ifu_io_imem_resp_valid; // @[Frontend.scala 106:20]
  wire [63:0] ifu_io_imem_resp_bits_rdata; // @[Frontend.scala 106:20]
  wire [81:0] ifu_io_imem_resp_bits_user; // @[Frontend.scala 106:20]
  wire  ifu_io_out_ready; // @[Frontend.scala 106:20]
  wire  ifu_io_out_valid; // @[Frontend.scala 106:20]
  wire [63:0] ifu_io_out_bits_instr; // @[Frontend.scala 106:20]
  wire [38:0] ifu_io_out_bits_pc; // @[Frontend.scala 106:20]
  wire [38:0] ifu_io_out_bits_pnpc; // @[Frontend.scala 106:20]
  wire  ifu_io_out_bits_exceptionVec_12; // @[Frontend.scala 106:20]
  wire [3:0] ifu_io_out_bits_brIdx; // @[Frontend.scala 106:20]
  wire [38:0] ifu_io_redirect_target; // @[Frontend.scala 106:20]
  wire  ifu_io_redirect_valid; // @[Frontend.scala 106:20]
  wire [3:0] ifu_io_flushVec; // @[Frontend.scala 106:20]
  wire  ifu_io_ipf; // @[Frontend.scala 106:20]
  wire  ifu_flushICache; // @[Frontend.scala 106:20]
  wire  ifu__T_243_valid; // @[Frontend.scala 106:20]
  wire [38:0] ifu__T_243_pc; // @[Frontend.scala 106:20]
  wire  ifu__T_243_isMissPredict; // @[Frontend.scala 106:20]
  wire [38:0] ifu__T_243_actualTarget; // @[Frontend.scala 106:20]
  wire  ifu__T_243_actualTaken; // @[Frontend.scala 106:20]
  wire [6:0] ifu__T_243_fuOpType; // @[Frontend.scala 106:20]
  wire [1:0] ifu__T_243_btbType; // @[Frontend.scala 106:20]
  wire  ifu__T_243_isRVC; // @[Frontend.scala 106:20]
  wire  ifu_DISPLAY_ENABLE; // @[Frontend.scala 106:20]
  wire  ifu__T_65_0; // @[Frontend.scala 106:20]
  wire  ifu_flushTLB; // @[Frontend.scala 106:20]
  wire  ifu__T_66_0; // @[Frontend.scala 106:20]
  wire  ibf_clock; // @[Frontend.scala 107:19]
  wire  ibf_reset; // @[Frontend.scala 107:19]
  wire  ibf_io_in_ready; // @[Frontend.scala 107:19]
  wire  ibf_io_in_valid; // @[Frontend.scala 107:19]
  wire [63:0] ibf_io_in_bits_instr; // @[Frontend.scala 107:19]
  wire [38:0] ibf_io_in_bits_pc; // @[Frontend.scala 107:19]
  wire [38:0] ibf_io_in_bits_pnpc; // @[Frontend.scala 107:19]
  wire  ibf_io_in_bits_exceptionVec_12; // @[Frontend.scala 107:19]
  wire [3:0] ibf_io_in_bits_brIdx; // @[Frontend.scala 107:19]
  wire  ibf_io_out_ready; // @[Frontend.scala 107:19]
  wire  ibf_io_out_valid; // @[Frontend.scala 107:19]
  wire [63:0] ibf_io_out_bits_instr; // @[Frontend.scala 107:19]
  wire [38:0] ibf_io_out_bits_pc; // @[Frontend.scala 107:19]
  wire [38:0] ibf_io_out_bits_pnpc; // @[Frontend.scala 107:19]
  wire  ibf_io_out_bits_exceptionVec_12; // @[Frontend.scala 107:19]
  wire [3:0] ibf_io_out_bits_brIdx; // @[Frontend.scala 107:19]
  wire  ibf_io_out_bits_crossPageIPFFix; // @[Frontend.scala 107:19]
  wire  ibf_io_flush; // @[Frontend.scala 107:19]
  wire  ibf_DISPLAY_ENABLE; // @[Frontend.scala 107:19]
  wire  idu_clock; // @[Frontend.scala 108:20]
  wire  idu_reset; // @[Frontend.scala 108:20]
  wire  idu_io_in_0_ready; // @[Frontend.scala 108:20]
  wire  idu_io_in_0_valid; // @[Frontend.scala 108:20]
  wire [63:0] idu_io_in_0_bits_instr; // @[Frontend.scala 108:20]
  wire [38:0] idu_io_in_0_bits_pc; // @[Frontend.scala 108:20]
  wire [38:0] idu_io_in_0_bits_pnpc; // @[Frontend.scala 108:20]
  wire  idu_io_in_0_bits_exceptionVec_12; // @[Frontend.scala 108:20]
  wire [3:0] idu_io_in_0_bits_brIdx; // @[Frontend.scala 108:20]
  wire  idu_io_in_0_bits_crossPageIPFFix; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_ready; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_valid; // @[Frontend.scala 108:20]
  wire [63:0] idu_io_out_0_bits_cf_instr; // @[Frontend.scala 108:20]
  wire [38:0] idu_io_out_0_bits_cf_pc; // @[Frontend.scala 108:20]
  wire [38:0] idu_io_out_0_bits_cf_pnpc; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_exceptionVec_1; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_exceptionVec_2; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_exceptionVec_12; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_0; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_1; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_2; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_3; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_4; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_5; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_6; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_7; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_8; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_9; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_10; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_11; // @[Frontend.scala 108:20]
  wire [3:0] idu_io_out_0_bits_cf_brIdx; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_crossPageIPFFix; // @[Frontend.scala 108:20]
  wire [1:0] idu_io_out_0_bits_ctrl_src1Type; // @[Frontend.scala 108:20]
  wire [1:0] idu_io_out_0_bits_ctrl_src2Type; // @[Frontend.scala 108:20]
  wire [2:0] idu_io_out_0_bits_ctrl_fuType; // @[Frontend.scala 108:20]
  wire [6:0] idu_io_out_0_bits_ctrl_fuOpType; // @[Frontend.scala 108:20]
  wire [4:0] idu_io_out_0_bits_ctrl_rfSrc1; // @[Frontend.scala 108:20]
  wire [4:0] idu_io_out_0_bits_ctrl_rfSrc2; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_ctrl_rfWen; // @[Frontend.scala 108:20]
  wire [4:0] idu_io_out_0_bits_ctrl_rfDest; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_ctrl_isNutCoreTrap; // @[Frontend.scala 108:20]
  wire [63:0] idu_io_out_0_bits_data_imm; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_0; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_1; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_2; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_3; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_4; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_5; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_6; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_7; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_8; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_9; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_10; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_11; // @[Frontend.scala 108:20]
  wire  idu__T_13; // @[Frontend.scala 108:20]
  wire  idu_vmEnable; // @[Frontend.scala 108:20]
  wire [11:0] idu_intrVec; // @[Frontend.scala 108:20]
  wire  idu__T_0; // @[Frontend.scala 108:20]
  wire  FlushableQueue_clock; // @[FlushableQueue.scala 104:21]
  wire  FlushableQueue_reset; // @[FlushableQueue.scala 104:21]
  wire  FlushableQueue_io_enq_ready; // @[FlushableQueue.scala 104:21]
  wire  FlushableQueue_io_enq_valid; // @[FlushableQueue.scala 104:21]
  wire [63:0] FlushableQueue_io_enq_bits_instr; // @[FlushableQueue.scala 104:21]
  wire [38:0] FlushableQueue_io_enq_bits_pc; // @[FlushableQueue.scala 104:21]
  wire [38:0] FlushableQueue_io_enq_bits_pnpc; // @[FlushableQueue.scala 104:21]
  wire  FlushableQueue_io_enq_bits_exceptionVec_12; // @[FlushableQueue.scala 104:21]
  wire [3:0] FlushableQueue_io_enq_bits_brIdx; // @[FlushableQueue.scala 104:21]
  wire  FlushableQueue_io_deq_ready; // @[FlushableQueue.scala 104:21]
  wire  FlushableQueue_io_deq_valid; // @[FlushableQueue.scala 104:21]
  wire [63:0] FlushableQueue_io_deq_bits_instr; // @[FlushableQueue.scala 104:21]
  wire [38:0] FlushableQueue_io_deq_bits_pc; // @[FlushableQueue.scala 104:21]
  wire [38:0] FlushableQueue_io_deq_bits_pnpc; // @[FlushableQueue.scala 104:21]
  wire  FlushableQueue_io_deq_bits_exceptionVec_12; // @[FlushableQueue.scala 104:21]
  wire [3:0] FlushableQueue_io_deq_bits_brIdx; // @[FlushableQueue.scala 104:21]
  wire  FlushableQueue_io_flush; // @[FlushableQueue.scala 104:21]
  wire  _T_1 = idu_io_out_0_ready & idu_io_out_0_valid; // @[Decoupled.scala 40:37]
  reg  _T_3; // @[Pipeline.scala 24:24]
  wire  _GEN_0 = _T_1 ? 1'h0 : _T_3; // @[Pipeline.scala 25:25]
  wire  _T_4 = ibf_io_out_valid & idu_io_in_0_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_1 = _T_4 | _GEN_0; // @[Pipeline.scala 26:38]
  reg [63:0] _T_6_instr; // @[Reg.scala 15:16]
  reg [38:0] _T_6_pc; // @[Reg.scala 15:16]
  reg [38:0] _T_6_pnpc; // @[Reg.scala 15:16]
  reg  _T_6_exceptionVec_12; // @[Reg.scala 15:16]
  reg [3:0] _T_6_brIdx; // @[Reg.scala 15:16]
  reg  _T_6_crossPageIPFFix; // @[Reg.scala 15:16]
  reg [63:0] _T_8; // @[GTimer.scala 24:20]
  wire [63:0] _T_10 = _T_8 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_14 = ~reset; // @[Debug.scala 56:24]
  reg [63:0] _T_17; // @[GTimer.scala 24:20]
  wire [63:0] _T_19 = _T_17 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_26; // @[GTimer.scala 24:20]
  wire [63:0] _T_28 = _T_26 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_30 = ifu_io_out_valid & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  reg [63:0] _T_35; // @[GTimer.scala 24:20]
  wire [63:0] _T_37 = _T_35 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_39 = idu_io_in_0_valid & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  IFU_inorder ifu ( // @[Frontend.scala 106:20]
    .clock(ifu_clock),
    .reset(ifu_reset),
    .io_imem_req_ready(ifu_io_imem_req_ready),
    .io_imem_req_valid(ifu_io_imem_req_valid),
    .io_imem_req_bits_addr(ifu_io_imem_req_bits_addr),
    .io_imem_req_bits_user(ifu_io_imem_req_bits_user),
    .io_imem_resp_ready(ifu_io_imem_resp_ready),
    .io_imem_resp_valid(ifu_io_imem_resp_valid),
    .io_imem_resp_bits_rdata(ifu_io_imem_resp_bits_rdata),
    .io_imem_resp_bits_user(ifu_io_imem_resp_bits_user),
    .io_out_ready(ifu_io_out_ready),
    .io_out_valid(ifu_io_out_valid),
    .io_out_bits_instr(ifu_io_out_bits_instr),
    .io_out_bits_pc(ifu_io_out_bits_pc),
    .io_out_bits_pnpc(ifu_io_out_bits_pnpc),
    .io_out_bits_exceptionVec_12(ifu_io_out_bits_exceptionVec_12),
    .io_out_bits_brIdx(ifu_io_out_bits_brIdx),
    .io_redirect_target(ifu_io_redirect_target),
    .io_redirect_valid(ifu_io_redirect_valid),
    .io_flushVec(ifu_io_flushVec),
    .io_ipf(ifu_io_ipf),
    .flushICache(ifu_flushICache),
    ._T_243_valid(ifu__T_243_valid),
    ._T_243_pc(ifu__T_243_pc),
    ._T_243_isMissPredict(ifu__T_243_isMissPredict),
    ._T_243_actualTarget(ifu__T_243_actualTarget),
    ._T_243_actualTaken(ifu__T_243_actualTaken),
    ._T_243_fuOpType(ifu__T_243_fuOpType),
    ._T_243_btbType(ifu__T_243_btbType),
    ._T_243_isRVC(ifu__T_243_isRVC),
    .DISPLAY_ENABLE(ifu_DISPLAY_ENABLE),
    ._T_65_0(ifu__T_65_0),
    .flushTLB(ifu_flushTLB),
    ._T_66_0(ifu__T_66_0)
  );
  NaiveRVCAlignBuffer ibf ( // @[Frontend.scala 107:19]
    .clock(ibf_clock),
    .reset(ibf_reset),
    .io_in_ready(ibf_io_in_ready),
    .io_in_valid(ibf_io_in_valid),
    .io_in_bits_instr(ibf_io_in_bits_instr),
    .io_in_bits_pc(ibf_io_in_bits_pc),
    .io_in_bits_pnpc(ibf_io_in_bits_pnpc),
    .io_in_bits_exceptionVec_12(ibf_io_in_bits_exceptionVec_12),
    .io_in_bits_brIdx(ibf_io_in_bits_brIdx),
    .io_out_ready(ibf_io_out_ready),
    .io_out_valid(ibf_io_out_valid),
    .io_out_bits_instr(ibf_io_out_bits_instr),
    .io_out_bits_pc(ibf_io_out_bits_pc),
    .io_out_bits_pnpc(ibf_io_out_bits_pnpc),
    .io_out_bits_exceptionVec_12(ibf_io_out_bits_exceptionVec_12),
    .io_out_bits_brIdx(ibf_io_out_bits_brIdx),
    .io_out_bits_crossPageIPFFix(ibf_io_out_bits_crossPageIPFFix),
    .io_flush(ibf_io_flush),
    .DISPLAY_ENABLE(ibf_DISPLAY_ENABLE)
  );
  IDU idu ( // @[Frontend.scala 108:20]
    .clock(idu_clock),
    .reset(idu_reset),
    .io_in_0_ready(idu_io_in_0_ready),
    .io_in_0_valid(idu_io_in_0_valid),
    .io_in_0_bits_instr(idu_io_in_0_bits_instr),
    .io_in_0_bits_pc(idu_io_in_0_bits_pc),
    .io_in_0_bits_pnpc(idu_io_in_0_bits_pnpc),
    .io_in_0_bits_exceptionVec_12(idu_io_in_0_bits_exceptionVec_12),
    .io_in_0_bits_brIdx(idu_io_in_0_bits_brIdx),
    .io_in_0_bits_crossPageIPFFix(idu_io_in_0_bits_crossPageIPFFix),
    .io_out_0_ready(idu_io_out_0_ready),
    .io_out_0_valid(idu_io_out_0_valid),
    .io_out_0_bits_cf_instr(idu_io_out_0_bits_cf_instr),
    .io_out_0_bits_cf_pc(idu_io_out_0_bits_cf_pc),
    .io_out_0_bits_cf_pnpc(idu_io_out_0_bits_cf_pnpc),
    .io_out_0_bits_cf_exceptionVec_1(idu_io_out_0_bits_cf_exceptionVec_1),
    .io_out_0_bits_cf_exceptionVec_2(idu_io_out_0_bits_cf_exceptionVec_2),
    .io_out_0_bits_cf_exceptionVec_12(idu_io_out_0_bits_cf_exceptionVec_12),
    .io_out_0_bits_cf_intrVec_0(idu_io_out_0_bits_cf_intrVec_0),
    .io_out_0_bits_cf_intrVec_1(idu_io_out_0_bits_cf_intrVec_1),
    .io_out_0_bits_cf_intrVec_2(idu_io_out_0_bits_cf_intrVec_2),
    .io_out_0_bits_cf_intrVec_3(idu_io_out_0_bits_cf_intrVec_3),
    .io_out_0_bits_cf_intrVec_4(idu_io_out_0_bits_cf_intrVec_4),
    .io_out_0_bits_cf_intrVec_5(idu_io_out_0_bits_cf_intrVec_5),
    .io_out_0_bits_cf_intrVec_6(idu_io_out_0_bits_cf_intrVec_6),
    .io_out_0_bits_cf_intrVec_7(idu_io_out_0_bits_cf_intrVec_7),
    .io_out_0_bits_cf_intrVec_8(idu_io_out_0_bits_cf_intrVec_8),
    .io_out_0_bits_cf_intrVec_9(idu_io_out_0_bits_cf_intrVec_9),
    .io_out_0_bits_cf_intrVec_10(idu_io_out_0_bits_cf_intrVec_10),
    .io_out_0_bits_cf_intrVec_11(idu_io_out_0_bits_cf_intrVec_11),
    .io_out_0_bits_cf_brIdx(idu_io_out_0_bits_cf_brIdx),
    .io_out_0_bits_cf_crossPageIPFFix(idu_io_out_0_bits_cf_crossPageIPFFix),
    .io_out_0_bits_ctrl_src1Type(idu_io_out_0_bits_ctrl_src1Type),
    .io_out_0_bits_ctrl_src2Type(idu_io_out_0_bits_ctrl_src2Type),
    .io_out_0_bits_ctrl_fuType(idu_io_out_0_bits_ctrl_fuType),
    .io_out_0_bits_ctrl_fuOpType(idu_io_out_0_bits_ctrl_fuOpType),
    .io_out_0_bits_ctrl_rfSrc1(idu_io_out_0_bits_ctrl_rfSrc1),
    .io_out_0_bits_ctrl_rfSrc2(idu_io_out_0_bits_ctrl_rfSrc2),
    .io_out_0_bits_ctrl_rfWen(idu_io_out_0_bits_ctrl_rfWen),
    .io_out_0_bits_ctrl_rfDest(idu_io_out_0_bits_ctrl_rfDest),
    .io_out_0_bits_ctrl_isNutCoreTrap(idu_io_out_0_bits_ctrl_isNutCoreTrap),
    .io_out_0_bits_data_imm(idu_io_out_0_bits_data_imm),
    .io_out_1_bits_cf_intrVec_0(idu_io_out_1_bits_cf_intrVec_0),
    .io_out_1_bits_cf_intrVec_1(idu_io_out_1_bits_cf_intrVec_1),
    .io_out_1_bits_cf_intrVec_2(idu_io_out_1_bits_cf_intrVec_2),
    .io_out_1_bits_cf_intrVec_3(idu_io_out_1_bits_cf_intrVec_3),
    .io_out_1_bits_cf_intrVec_4(idu_io_out_1_bits_cf_intrVec_4),
    .io_out_1_bits_cf_intrVec_5(idu_io_out_1_bits_cf_intrVec_5),
    .io_out_1_bits_cf_intrVec_6(idu_io_out_1_bits_cf_intrVec_6),
    .io_out_1_bits_cf_intrVec_7(idu_io_out_1_bits_cf_intrVec_7),
    .io_out_1_bits_cf_intrVec_8(idu_io_out_1_bits_cf_intrVec_8),
    .io_out_1_bits_cf_intrVec_9(idu_io_out_1_bits_cf_intrVec_9),
    .io_out_1_bits_cf_intrVec_10(idu_io_out_1_bits_cf_intrVec_10),
    .io_out_1_bits_cf_intrVec_11(idu_io_out_1_bits_cf_intrVec_11),
    ._T_13(idu__T_13),
    .vmEnable(idu_vmEnable),
    .intrVec(idu_intrVec),
    ._T_0(idu__T_0)
  );
  FlushableQueue FlushableQueue ( // @[FlushableQueue.scala 104:21]
    .clock(FlushableQueue_clock),
    .reset(FlushableQueue_reset),
    .io_enq_ready(FlushableQueue_io_enq_ready),
    .io_enq_valid(FlushableQueue_io_enq_valid),
    .io_enq_bits_instr(FlushableQueue_io_enq_bits_instr),
    .io_enq_bits_pc(FlushableQueue_io_enq_bits_pc),
    .io_enq_bits_pnpc(FlushableQueue_io_enq_bits_pnpc),
    .io_enq_bits_exceptionVec_12(FlushableQueue_io_enq_bits_exceptionVec_12),
    .io_enq_bits_brIdx(FlushableQueue_io_enq_bits_brIdx),
    .io_deq_ready(FlushableQueue_io_deq_ready),
    .io_deq_valid(FlushableQueue_io_deq_valid),
    .io_deq_bits_instr(FlushableQueue_io_deq_bits_instr),
    .io_deq_bits_pc(FlushableQueue_io_deq_bits_pc),
    .io_deq_bits_pnpc(FlushableQueue_io_deq_bits_pnpc),
    .io_deq_bits_exceptionVec_12(FlushableQueue_io_deq_bits_exceptionVec_12),
    .io_deq_bits_brIdx(FlushableQueue_io_deq_bits_brIdx),
    .io_flush(FlushableQueue_io_flush)
  );
  assign io_out_0_valid = idu_io_out_0_valid; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_instr = idu_io_out_0_bits_cf_instr; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_pc = idu_io_out_0_bits_cf_pc; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_pnpc = idu_io_out_0_bits_cf_pnpc; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_exceptionVec_1 = idu_io_out_0_bits_cf_exceptionVec_1; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_exceptionVec_2 = idu_io_out_0_bits_cf_exceptionVec_2; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_exceptionVec_12 = idu_io_out_0_bits_cf_exceptionVec_12; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_0 = idu_io_out_0_bits_cf_intrVec_0; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_1 = idu_io_out_0_bits_cf_intrVec_1; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_2 = idu_io_out_0_bits_cf_intrVec_2; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_3 = idu_io_out_0_bits_cf_intrVec_3; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_4 = idu_io_out_0_bits_cf_intrVec_4; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_5 = idu_io_out_0_bits_cf_intrVec_5; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_6 = idu_io_out_0_bits_cf_intrVec_6; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_7 = idu_io_out_0_bits_cf_intrVec_7; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_8 = idu_io_out_0_bits_cf_intrVec_8; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_9 = idu_io_out_0_bits_cf_intrVec_9; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_10 = idu_io_out_0_bits_cf_intrVec_10; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_11 = idu_io_out_0_bits_cf_intrVec_11; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_brIdx = idu_io_out_0_bits_cf_brIdx; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_crossPageIPFFix = idu_io_out_0_bits_cf_crossPageIPFFix; // @[Frontend.scala 120:10]
  assign io_out_0_bits_ctrl_src1Type = idu_io_out_0_bits_ctrl_src1Type; // @[Frontend.scala 120:10]
  assign io_out_0_bits_ctrl_src2Type = idu_io_out_0_bits_ctrl_src2Type; // @[Frontend.scala 120:10]
  assign io_out_0_bits_ctrl_fuType = idu_io_out_0_bits_ctrl_fuType; // @[Frontend.scala 120:10]
  assign io_out_0_bits_ctrl_fuOpType = idu_io_out_0_bits_ctrl_fuOpType; // @[Frontend.scala 120:10]
  assign io_out_0_bits_ctrl_rfSrc1 = idu_io_out_0_bits_ctrl_rfSrc1; // @[Frontend.scala 120:10]
  assign io_out_0_bits_ctrl_rfSrc2 = idu_io_out_0_bits_ctrl_rfSrc2; // @[Frontend.scala 120:10]
  assign io_out_0_bits_ctrl_rfWen = idu_io_out_0_bits_ctrl_rfWen; // @[Frontend.scala 120:10]
  assign io_out_0_bits_ctrl_rfDest = idu_io_out_0_bits_ctrl_rfDest; // @[Frontend.scala 120:10]
  assign io_out_0_bits_ctrl_isNutCoreTrap = idu_io_out_0_bits_ctrl_isNutCoreTrap; // @[Frontend.scala 120:10]
  assign io_out_0_bits_data_imm = idu_io_out_0_bits_data_imm; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_0 = idu_io_out_1_bits_cf_intrVec_0; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_1 = idu_io_out_1_bits_cf_intrVec_1; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_2 = idu_io_out_1_bits_cf_intrVec_2; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_3 = idu_io_out_1_bits_cf_intrVec_3; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_4 = idu_io_out_1_bits_cf_intrVec_4; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_5 = idu_io_out_1_bits_cf_intrVec_5; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_6 = idu_io_out_1_bits_cf_intrVec_6; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_7 = idu_io_out_1_bits_cf_intrVec_7; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_8 = idu_io_out_1_bits_cf_intrVec_8; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_9 = idu_io_out_1_bits_cf_intrVec_9; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_10 = idu_io_out_1_bits_cf_intrVec_10; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_11 = idu_io_out_1_bits_cf_intrVec_11; // @[Frontend.scala 120:10]
  assign io_imem_req_valid = ifu_io_imem_req_valid; // @[Frontend.scala 125:11]
  assign io_imem_req_bits_addr = ifu_io_imem_req_bits_addr; // @[Frontend.scala 125:11]
  assign io_imem_req_bits_user = {{5'd0}, ifu_io_imem_req_bits_user}; // @[Frontend.scala 125:11]
  assign io_imem_resp_ready = ifu_io_imem_resp_ready; // @[Frontend.scala 125:11]
  assign io_flushVec = ifu_io_flushVec; // @[Frontend.scala 122:15]
  assign _T_0 = idu__T_0;
  assign _T_65 = ifu__T_65_0;
  assign _T_66 = ifu__T_66_0;
  assign ifu_clock = clock;
  assign ifu_reset = reset;
  assign ifu_io_imem_req_ready = io_imem_req_ready; // @[Frontend.scala 125:11]
  assign ifu_io_imem_resp_valid = io_imem_resp_valid; // @[Frontend.scala 125:11]
  assign ifu_io_imem_resp_bits_rdata = io_imem_resp_bits_rdata; // @[Frontend.scala 125:11]
  assign ifu_io_imem_resp_bits_user = io_imem_resp_bits_user[81:0]; // @[Frontend.scala 125:11]
  assign ifu_io_out_ready = FlushableQueue_io_enq_ready; // @[FlushableQueue.scala 108:17]
  assign ifu_io_redirect_target = io_redirect_target; // @[Frontend.scala 121:15]
  assign ifu_io_redirect_valid = io_redirect_valid; // @[Frontend.scala 121:15]
  assign ifu_io_ipf = io_ipf; // @[Frontend.scala 124:10]
  assign ifu_flushICache = flushICache;
  assign ifu__T_243_valid = _T_243_valid;
  assign ifu__T_243_pc = _T_243_pc;
  assign ifu__T_243_isMissPredict = _T_243_isMissPredict;
  assign ifu__T_243_actualTarget = _T_243_actualTarget;
  assign ifu__T_243_actualTaken = _T_243_actualTaken;
  assign ifu__T_243_fuOpType = _T_243_fuOpType;
  assign ifu__T_243_btbType = _T_243_btbType;
  assign ifu__T_243_isRVC = _T_243_isRVC;
  assign ifu_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign ifu_flushTLB = flushTLB;
  assign ibf_clock = clock;
  assign ibf_reset = reset;
  assign ibf_io_in_valid = FlushableQueue_io_deq_valid; // @[Frontend.scala 112:11]
  assign ibf_io_in_bits_instr = FlushableQueue_io_deq_bits_instr; // @[Frontend.scala 112:11]
  assign ibf_io_in_bits_pc = FlushableQueue_io_deq_bits_pc; // @[Frontend.scala 112:11]
  assign ibf_io_in_bits_pnpc = FlushableQueue_io_deq_bits_pnpc; // @[Frontend.scala 112:11]
  assign ibf_io_in_bits_exceptionVec_12 = FlushableQueue_io_deq_bits_exceptionVec_12; // @[Frontend.scala 112:11]
  assign ibf_io_in_bits_brIdx = FlushableQueue_io_deq_bits_brIdx; // @[Frontend.scala 112:11]
  assign ibf_io_out_ready = idu_io_in_0_ready; // @[Pipeline.scala 29:16]
  assign ibf_io_flush = ifu_io_flushVec[1]; // @[Frontend.scala 119:16]
  assign ibf_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign idu_clock = clock;
  assign idu_reset = reset;
  assign idu_io_in_0_valid = _T_3; // @[Pipeline.scala 31:17]
  assign idu_io_in_0_bits_instr = _T_6_instr; // @[Pipeline.scala 30:16]
  assign idu_io_in_0_bits_pc = _T_6_pc; // @[Pipeline.scala 30:16]
  assign idu_io_in_0_bits_pnpc = _T_6_pnpc; // @[Pipeline.scala 30:16]
  assign idu_io_in_0_bits_exceptionVec_12 = _T_6_exceptionVec_12; // @[Pipeline.scala 30:16]
  assign idu_io_in_0_bits_brIdx = _T_6_brIdx; // @[Pipeline.scala 30:16]
  assign idu_io_in_0_bits_crossPageIPFFix = _T_6_crossPageIPFFix; // @[Pipeline.scala 30:16]
  assign idu_io_out_0_ready = io_out_0_ready; // @[Frontend.scala 120:10]
  assign idu__T_13 = DISPLAY_ENABLE;
  assign idu_vmEnable = vmEnable;
  assign idu_intrVec = intrVec;
  assign FlushableQueue_clock = clock;
  assign FlushableQueue_reset = reset;
  assign FlushableQueue_io_enq_valid = ifu_io_out_valid; // @[FlushableQueue.scala 105:22]
  assign FlushableQueue_io_enq_bits_instr = ifu_io_out_bits_instr; // @[FlushableQueue.scala 106:21]
  assign FlushableQueue_io_enq_bits_pc = ifu_io_out_bits_pc; // @[FlushableQueue.scala 106:21]
  assign FlushableQueue_io_enq_bits_pnpc = ifu_io_out_bits_pnpc; // @[FlushableQueue.scala 106:21]
  assign FlushableQueue_io_enq_bits_exceptionVec_12 = ifu_io_out_bits_exceptionVec_12; // @[FlushableQueue.scala 106:21]
  assign FlushableQueue_io_enq_bits_brIdx = ifu_io_out_bits_brIdx; // @[FlushableQueue.scala 106:21]
  assign FlushableQueue_io_deq_ready = ibf_io_in_ready; // @[Frontend.scala 112:11]
  assign FlushableQueue_io_flush = ifu_io_flushVec[0]; // @[FlushableQueue.scala 107:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_3 = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  _T_6_instr = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  _T_6_pc = _RAND_2[38:0];
  _RAND_3 = {2{`RANDOM}};
  _T_6_pnpc = _RAND_3[38:0];
  _RAND_4 = {1{`RANDOM}};
  _T_6_exceptionVec_12 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _T_6_brIdx = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  _T_6_crossPageIPFFix = _RAND_6[0:0];
  _RAND_7 = {2{`RANDOM}};
  _T_8 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  _T_17 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  _T_26 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  _T_35 = _RAND_10[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_3 <= 1'h0;
    end else if (ifu_io_flushVec[1]) begin
      _T_3 <= 1'h0;
    end else begin
      _T_3 <= _GEN_1;
    end
    if (_T_4) begin
      _T_6_instr <= ibf_io_out_bits_instr;
    end
    if (_T_4) begin
      _T_6_pc <= ibf_io_out_bits_pc;
    end
    if (_T_4) begin
      _T_6_pnpc <= ibf_io_out_bits_pnpc;
    end
    if (_T_4) begin
      _T_6_exceptionVec_12 <= ibf_io_out_bits_exceptionVec_12;
    end
    if (_T_4) begin
      _T_6_brIdx <= ibf_io_out_bits_brIdx;
    end
    if (_T_4) begin
      _T_6_crossPageIPFFix <= ibf_io_out_bits_crossPageIPFFix;
    end
    if (reset) begin
      _T_8 <= 64'h0;
    end else begin
      _T_8 <= _T_10;
    end
    if (reset) begin
      _T_17 <= 64'h0;
    end else begin
      _T_17 <= _T_19;
    end
    if (reset) begin
      _T_26 <= 64'h0;
    end else begin
      _T_26 <= _T_28;
    end
    if (reset) begin
      _T_35 <= 64'h0;
    end else begin
      _T_35 <= _T_37;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_14) begin
          $fwrite(32'h80000002,"[%d] Frontend_inorder: ",_T_8); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_14) begin
          $fwrite(32'h80000002,"------------------------ FRONTEND:------------------------\n"); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_14) begin
          $fwrite(32'h80000002,"[%d] Frontend_inorder: ",_T_17); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_14) begin
          $fwrite(32'h80000002,"flush = %b, ifu:(%d,%d), idu:(%d,%d)\n",ifu_io_flushVec,ifu_io_out_valid,ifu_io_out_ready,idu_io_in_0_valid,idu_io_in_0_ready); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_30 & _T_14) begin
          $fwrite(32'h80000002,"[%d] Frontend_inorder: ",_T_26); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_30 & _T_14) begin
          $fwrite(32'h80000002,"IFU: pc = 0x%x, instr = 0x%x\n",ifu_io_out_bits_pc,ifu_io_out_bits_instr); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & _T_14) begin
          $fwrite(32'h80000002,"[%d] Frontend_inorder: ",_T_35); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_39 & _T_14) begin
          $fwrite(32'h80000002,"IDU1: pc = 0x%x, instr = 0x%x, pnpc = 0x%x\n",idu_io_in_0_bits_pc,idu_io_in_0_bits_instr,idu_io_in_0_bits_pnpc); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ISU(
  input         clock,
  input         reset,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [63:0] io_in_0_bits_cf_instr,
  input  [38:0] io_in_0_bits_cf_pc,
  input  [38:0] io_in_0_bits_cf_pnpc,
  input         io_in_0_bits_cf_exceptionVec_1,
  input         io_in_0_bits_cf_exceptionVec_2,
  input         io_in_0_bits_cf_exceptionVec_12,
  input         io_in_0_bits_cf_intrVec_0,
  input         io_in_0_bits_cf_intrVec_1,
  input         io_in_0_bits_cf_intrVec_2,
  input         io_in_0_bits_cf_intrVec_3,
  input         io_in_0_bits_cf_intrVec_4,
  input         io_in_0_bits_cf_intrVec_5,
  input         io_in_0_bits_cf_intrVec_6,
  input         io_in_0_bits_cf_intrVec_7,
  input         io_in_0_bits_cf_intrVec_8,
  input         io_in_0_bits_cf_intrVec_9,
  input         io_in_0_bits_cf_intrVec_10,
  input         io_in_0_bits_cf_intrVec_11,
  input  [3:0]  io_in_0_bits_cf_brIdx,
  input         io_in_0_bits_cf_crossPageIPFFix,
  input  [1:0]  io_in_0_bits_ctrl_src1Type,
  input  [1:0]  io_in_0_bits_ctrl_src2Type,
  input  [2:0]  io_in_0_bits_ctrl_fuType,
  input  [6:0]  io_in_0_bits_ctrl_fuOpType,
  input  [4:0]  io_in_0_bits_ctrl_rfSrc1,
  input  [4:0]  io_in_0_bits_ctrl_rfSrc2,
  input         io_in_0_bits_ctrl_rfWen,
  input  [4:0]  io_in_0_bits_ctrl_rfDest,
  input         io_in_0_bits_ctrl_isNutCoreTrap,
  input  [63:0] io_in_0_bits_data_imm,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_cf_instr,
  output [38:0] io_out_bits_cf_pc,
  output [38:0] io_out_bits_cf_pnpc,
  output        io_out_bits_cf_exceptionVec_1,
  output        io_out_bits_cf_exceptionVec_2,
  output        io_out_bits_cf_exceptionVec_12,
  output        io_out_bits_cf_intrVec_0,
  output        io_out_bits_cf_intrVec_1,
  output        io_out_bits_cf_intrVec_2,
  output        io_out_bits_cf_intrVec_3,
  output        io_out_bits_cf_intrVec_4,
  output        io_out_bits_cf_intrVec_5,
  output        io_out_bits_cf_intrVec_6,
  output        io_out_bits_cf_intrVec_7,
  output        io_out_bits_cf_intrVec_8,
  output        io_out_bits_cf_intrVec_9,
  output        io_out_bits_cf_intrVec_10,
  output        io_out_bits_cf_intrVec_11,
  output [3:0]  io_out_bits_cf_brIdx,
  output        io_out_bits_cf_crossPageIPFFix,
  output [2:0]  io_out_bits_ctrl_fuType,
  output [6:0]  io_out_bits_ctrl_fuOpType,
  output        io_out_bits_ctrl_rfWen,
  output [4:0]  io_out_bits_ctrl_rfDest,
  output        io_out_bits_ctrl_isNutCoreTrap,
  output [63:0] io_out_bits_data_src1,
  output [63:0] io_out_bits_data_src2,
  output [63:0] io_out_bits_data_imm,
  output [63:0] io_out_bits_data_srf_0,
  output [63:0] io_out_bits_data_srf_1,
  output [63:0] io_out_bits_data_srf_2,
  output [63:0] io_out_bits_data_srf_3,
  input         io_wb_rfWen,
  input  [4:0]  io_wb_rfDest,
  input  [63:0] io_wb_rfData,
  input         io_wb_srfWen,
  input  [2:0]  io_wb_srfDest,
  input  [63:0] io_wb_srfData,
  input         io_forward_valid,
  input         io_forward_wb_rfWen,
  input  [4:0]  io_forward_wb_rfDest,
  input  [63:0] io_forward_wb_rfData,
  input  [2:0]  io_forward_wb_srfDest,
  input  [63:0] io_forward_wb_srfData,
  input  [2:0]  io_forward_fuType,
  input         io_flush,
  output        _T_183_0,
  output [63:0] _T_284_0_0,
  output [63:0] _T_284_0_1,
  output [63:0] _T_284_0_2,
  output [63:0] _T_284_0_3,
  output [63:0] _T_284_0_4,
  output [63:0] _T_284_0_5,
  output [63:0] _T_284_0_6,
  output [63:0] _T_284_0_7,
  output [63:0] _T_284_0_8,
  output [63:0] _T_284_0_9,
  output [63:0] _T_284_0_10,
  output [63:0] _T_284_0_11,
  output [63:0] _T_284_0_12,
  output [63:0] _T_284_0_13,
  output [63:0] _T_284_0_14,
  output [63:0] _T_284_0_15,
  output [63:0] _T_284_0_16,
  output [63:0] _T_284_0_17,
  output [63:0] _T_284_0_18,
  output [63:0] _T_284_0_19,
  output [63:0] _T_284_0_20,
  output [63:0] _T_284_0_21,
  output [63:0] _T_284_0_22,
  output [63:0] _T_284_0_23,
  output [63:0] _T_284_0_24,
  output [63:0] _T_284_0_25,
  output [63:0] _T_284_0_26,
  output [63:0] _T_284_0_27,
  output [63:0] _T_284_0_28,
  output [63:0] _T_284_0_29,
  output [63:0] _T_284_0_30,
  output [63:0] _T_284_0_31,
  output        _T_186_0,
  input         DISPLAY_ENABLE,
  output        _T_187_0
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] _T_31 [0:31]; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_84_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_84_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_103_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_103_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_189_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_189_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_192_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_192_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_195_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_195_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_198_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_198_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_201_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_201_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_204_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_204_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_207_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_207_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_210_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_210_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_213_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_213_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_216_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_216_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_219_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_219_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_222_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_222_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_225_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_225_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_228_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_228_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_231_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_231_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_234_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_234_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_237_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_237_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_240_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_240_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_243_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_243_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_246_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_246_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_249_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_249_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_252_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_252_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_255_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_255_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_258_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_258_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_261_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_261_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_264_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_264_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_267_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_267_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_270_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_270_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_273_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_273_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_276_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_276_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_279_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_279_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_282_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_282_addr; // @[RF.scala 31:15]
  wire [63:0] _T_31__T_113_data; // @[RF.scala 31:15]
  wire [4:0] _T_31__T_113_addr; // @[RF.scala 31:15]
  wire  _T_31__T_113_mask; // @[RF.scala 31:15]
  wire  _T_31__T_113_en; // @[RF.scala 31:15]
  reg [63:0] _T_32 [0:5]; // @[RF.scala 50:16]
  wire [63:0] _T_32__T_46_data; // @[RF.scala 50:16]
  wire [2:0] _T_32__T_46_addr; // @[RF.scala 50:16]
  wire [63:0] _T_32__T_51_data; // @[RF.scala 50:16]
  wire [2:0] _T_32__T_51_addr; // @[RF.scala 50:16]
  wire [63:0] _T_32__T_56_data; // @[RF.scala 50:16]
  wire [2:0] _T_32__T_56_addr; // @[RF.scala 50:16]
  wire [63:0] _T_32__T_61_data; // @[RF.scala 50:16]
  wire [2:0] _T_32__T_61_addr; // @[RF.scala 50:16]
  wire [63:0] _T_32__T_66_data; // @[RF.scala 50:16]
  wire [2:0] _T_32__T_66_addr; // @[RF.scala 50:16]
  wire [63:0] _T_32__T_118_data; // @[RF.scala 50:16]
  wire [2:0] _T_32__T_118_addr; // @[RF.scala 50:16]
  wire [63:0] _T_32__T_121_data; // @[RF.scala 50:16]
  wire [2:0] _T_32__T_121_addr; // @[RF.scala 50:16]
  wire [63:0] _T_32__T_124_data; // @[RF.scala 50:16]
  wire [2:0] _T_32__T_124_addr; // @[RF.scala 50:16]
  wire [63:0] _T_32__T_127_data; // @[RF.scala 50:16]
  wire [2:0] _T_32__T_127_addr; // @[RF.scala 50:16]
  wire [63:0] _T_32__T_130_data; // @[RF.scala 50:16]
  wire [2:0] _T_32__T_130_addr; // @[RF.scala 50:16]
  wire [63:0] _T_32__T_69_data; // @[RF.scala 50:16]
  wire [2:0] _T_32__T_69_addr; // @[RF.scala 50:16]
  wire  _T_32__T_69_mask; // @[RF.scala 50:16]
  wire  _T_32__T_69_en; // @[RF.scala 50:16]
  wire  forwardRfWen = io_forward_wb_rfWen & io_forward_valid; // @[ISU.scala 44:42]
  wire  _T = io_forward_fuType != 3'h0; // @[ISU.scala 45:41]
  wire  _T_1 = io_forward_fuType != 3'h1; // @[ISU.scala 45:79]
  wire  dontForward1 = _T & _T_1; // @[ISU.scala 45:57]
  wire  _T_2 = io_in_0_bits_ctrl_rfSrc1 != 5'h0; // @[ISU.scala 42:69]
  wire  _T_3 = io_in_0_bits_ctrl_rfSrc1 == io_forward_wb_rfDest; // @[ISU.scala 42:88]
  wire  _T_4 = _T_2 & _T_3; // @[ISU.scala 42:78]
  wire  src1DependEX = _T_4 & forwardRfWen; // @[ISU.scala 42:100]
  wire  _T_5 = io_in_0_bits_ctrl_rfSrc2 != 5'h0; // @[ISU.scala 42:69]
  wire  _T_6 = io_in_0_bits_ctrl_rfSrc2 == io_forward_wb_rfDest; // @[ISU.scala 42:88]
  wire  _T_7 = _T_5 & _T_6; // @[ISU.scala 42:78]
  wire  src2DependEX = _T_7 & forwardRfWen; // @[ISU.scala 42:100]
  wire  _T_9 = io_in_0_bits_ctrl_rfSrc1 == io_wb_rfDest; // @[ISU.scala 42:88]
  wire  _T_10 = _T_2 & _T_9; // @[ISU.scala 42:78]
  wire  src1DependWB = _T_10 & io_wb_rfWen; // @[ISU.scala 42:100]
  wire  _T_12 = io_in_0_bits_ctrl_rfSrc2 == io_wb_rfDest; // @[ISU.scala 42:88]
  wire  _T_13 = _T_5 & _T_12; // @[ISU.scala 42:78]
  wire  src2DependWB = _T_13 & io_wb_rfWen; // @[ISU.scala 42:100]
  wire  _T_14 = ~dontForward1; // @[ISU.scala 51:46]
  wire  src1ForwardNextCycle = src1DependEX & _T_14; // @[ISU.scala 51:43]
  wire  src2ForwardNextCycle = src2DependEX & _T_14; // @[ISU.scala 52:43]
  wire  _T_16 = ~src1DependEX; // @[ISU.scala 53:55]
  wire  _T_17 = dontForward1 ? _T_16 : 1'h1; // @[ISU.scala 53:40]
  wire  src1Forward = src1DependWB & _T_17; // @[ISU.scala 53:34]
  wire  _T_18 = ~src2DependEX; // @[ISU.scala 54:55]
  wire  _T_19 = dontForward1 ? _T_18 : 1'h1; // @[ISU.scala 54:40]
  wire  src2Forward = src2DependWB & _T_19; // @[ISU.scala 54:34]
  reg [31:0] _T_20; // @[RF.scala 37:21]
  wire [31:0] _T_21 = _T_20 >> io_in_0_bits_ctrl_rfSrc1; // @[RF.scala 38:37]
  wire  _T_23 = ~_T_21[0]; // @[ISU.scala 57:19]
  wire  _T_24 = _T_23 | src1ForwardNextCycle; // @[ISU.scala 57:38]
  wire  src1Ready = _T_24 | src1Forward; // @[ISU.scala 57:62]
  wire [31:0] _T_25 = _T_20 >> io_in_0_bits_ctrl_rfSrc2; // @[RF.scala 38:37]
  wire  _T_27 = ~_T_25[0]; // @[ISU.scala 58:19]
  wire  _T_28 = _T_27 | src2ForwardNextCycle; // @[ISU.scala 58:38]
  wire  src2Ready = _T_28 | src2Forward; // @[ISU.scala 58:62]
  wire  _T_29 = io_in_0_valid & src1Ready; // @[ISU.scala 59:34]
  wire  _T_33 = 7'h4 == io_in_0_bits_ctrl_fuOpType; // @[LookupTree.scala 24:34]
  wire  _T_34 = 7'h9 == io_in_0_bits_ctrl_fuOpType; // @[LookupTree.scala 24:34]
  wire  _T_35 = 7'h19 == io_in_0_bits_ctrl_fuOpType; // @[LookupTree.scala 24:34]
  wire  _T_36 = 7'h2 == io_in_0_bits_ctrl_fuOpType; // @[LookupTree.scala 24:34]
  wire [1:0] _T_38 = _T_34 ? 2'h3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_39 = _T_35 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_40 = _T_36 ? 3'h5 : 3'h0; // @[Mux.scala 27:72]
  wire [1:0] _GEN_23 = {{1'd0}, _T_33}; // @[Mux.scala 27:72]
  wire [1:0] _T_41 = _GEN_23 | _T_38; // @[Mux.scala 27:72]
  wire [1:0] _T_42 = _T_41 | _T_39; // @[Mux.scala 27:72]
  wire [2:0] _GEN_24 = {{1'd0}, _T_42}; // @[Mux.scala 27:72]
  wire [2:0] srfReq = _GEN_24 | _T_40; // @[Mux.scala 27:72]
  wire  _T_44 = io_forward_wb_srfDest == srfReq; // @[ISU.scala 71:66]
  wire  _T_45 = io_wb_srfDest == srfReq; // @[ISU.scala 72:63]
  wire [63:0] _T_47 = _T_45 ? io_wb_srfData : _T_32__T_46_data; // @[ISU.scala 72:48]
  wire [63:0] _T_52 = _T_45 ? io_wb_srfData : _T_32__T_51_data; // @[ISU.scala 74:48]
  wire [63:0] _T_57 = _T_45 ? io_wb_srfData : _T_32__T_56_data; // @[ISU.scala 76:48]
  wire [63:0] _T_67 = _T_45 ? io_wb_srfData : _T_32__T_66_data; // @[ISU.scala 80:48]
  wire  _T_71 = io_in_0_bits_ctrl_src1Type == 2'h1; // @[ISU.scala 85:34]
  wire [24:0] _T_74 = io_in_0_bits_cf_pc[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_75 = {_T_74,io_in_0_bits_cf_pc}; // @[Cat.scala 29:58]
  wire  _T_76 = ~src1ForwardNextCycle; // @[ISU.scala 87:21]
  wire  _T_77 = src1Forward & _T_76; // @[ISU.scala 87:18]
  wire  _T_78 = io_in_0_bits_ctrl_src1Type != 2'h1; // @[ISU.scala 88:35]
  wire  _T_80 = _T_78 & _T_76; // @[ISU.scala 88:51]
  wire  _T_81 = ~src1Forward; // @[ISU.scala 88:79]
  wire  _T_82 = _T_80 & _T_81; // @[ISU.scala 88:76]
  wire  _T_83 = io_in_0_bits_ctrl_rfSrc1 == 5'h0; // @[RF.scala 32:42]
  wire [63:0] _T_85 = _T_83 ? 64'h0 : _T_31__T_84_data; // @[RF.scala 32:36]
  wire [63:0] _T_86 = _T_71 ? _T_75 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_87 = src1ForwardNextCycle ? io_forward_wb_rfData : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_88 = _T_77 ? io_wb_rfData : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_89 = _T_82 ? _T_85 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_90 = _T_86 | _T_87; // @[Mux.scala 27:72]
  wire [63:0] _T_91 = _T_90 | _T_88; // @[Mux.scala 27:72]
  wire  _T_94 = io_in_0_bits_ctrl_src2Type != 2'h0; // @[ISU.scala 91:34]
  wire  _T_95 = ~src2ForwardNextCycle; // @[ISU.scala 93:21]
  wire  _T_96 = src2Forward & _T_95; // @[ISU.scala 93:18]
  wire  _T_97 = io_in_0_bits_ctrl_src2Type == 2'h0; // @[ISU.scala 94:35]
  wire  _T_99 = _T_97 & _T_95; // @[ISU.scala 94:52]
  wire  _T_100 = ~src2Forward; // @[ISU.scala 94:80]
  wire  _T_101 = _T_99 & _T_100; // @[ISU.scala 94:77]
  wire  _T_102 = io_in_0_bits_ctrl_rfSrc2 == 5'h0; // @[RF.scala 32:42]
  wire [63:0] _T_104 = _T_102 ? 64'h0 : _T_31__T_103_data; // @[RF.scala 32:36]
  wire [63:0] _T_105 = _T_94 ? io_in_0_bits_data_imm : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_106 = src2ForwardNextCycle ? io_forward_wb_rfData : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_107 = _T_96 ? io_wb_rfData : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_108 = _T_101 ? _T_104 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_109 = _T_105 | _T_106; // @[Mux.scala 27:72]
  wire [63:0] _T_110 = _T_109 | _T_107; // @[Mux.scala 27:72]
  wire  _T_120 = ~reset; // @[ISU.scala 113:13]
  wire  _T_147 = io_wb_rfDest != 5'h0; // @[ISU.scala 42:69]
  wire  _T_148 = io_wb_rfDest == io_forward_wb_rfDest; // @[ISU.scala 42:88]
  wire  _T_149 = _T_147 & _T_148; // @[ISU.scala 42:78]
  wire  _T_150 = _T_149 & forwardRfWen; // @[ISU.scala 42:100]
  wire  _T_151 = ~_T_150; // @[ISU.scala 127:40]
  wire  _T_152 = io_wb_rfWen & _T_151; // @[ISU.scala 127:37]
  wire [62:0] _T_153 = 63'h1 << io_wb_rfDest; // @[RF.scala 39:39]
  wire [31:0] wbClearMask = _T_152 ? _T_153[31:0] : 32'h0; // @[ISU.scala 127:24]
  wire  _T_155 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire [62:0] _T_156 = 63'h1 << io_in_0_bits_ctrl_rfDest; // @[RF.scala 39:39]
  wire [31:0] isuFireSetMask = _T_155 ? _T_156[31:0] : 32'h0; // @[ISU.scala 129:27]
  wire [31:0] _T_164 = ~wbClearMask; // @[RF.scala 45:26]
  wire [31:0] _T_165 = _T_20 & _T_164; // @[RF.scala 45:24]
  wire [31:0] _T_166 = _T_165 | isuFireSetMask; // @[RF.scala 45:38]
  wire [31:0] _T_168 = {_T_166[31:1],1'h0}; // @[Cat.scala 29:58]
  wire  _T_169 = ~io_in_0_valid; // @[ISU.scala 133:21]
  reg [63:0] _T_173; // @[GTimer.scala 24:20]
  wire [63:0] _T_175 = _T_173 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_177 = _T_155 & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  wire  _T_182 = ~io_out_valid; // @[ISU.scala 139:43]
  wire  _T_183 = io_in_0_valid & _T_182; // @[ISU.scala 139:40]
  wire  _T_185 = ~_T_155; // @[ISU.scala 140:41]
  wire  _T_186 = io_out_valid & _T_185; // @[ISU.scala 140:38]
  wire  _T_187 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire [63:0] _T_190 = 64'h0; // @[RF.scala 32:36]
  wire [63:0] _T_193 = _T_31__T_192_data; // @[RF.scala 32:36]
  wire [63:0] _T_196 = _T_31__T_195_data; // @[RF.scala 32:36]
  wire [63:0] _T_199 = _T_31__T_198_data; // @[RF.scala 32:36]
  wire [63:0] _T_202 = _T_31__T_201_data; // @[RF.scala 32:36]
  wire [63:0] _T_205 = _T_31__T_204_data; // @[RF.scala 32:36]
  wire [63:0] _T_208 = _T_31__T_207_data; // @[RF.scala 32:36]
  wire [63:0] _T_211 = _T_31__T_210_data; // @[RF.scala 32:36]
  wire [63:0] _T_214 = _T_31__T_213_data; // @[RF.scala 32:36]
  wire [63:0] _T_217 = _T_31__T_216_data; // @[RF.scala 32:36]
  wire [63:0] _T_220 = _T_31__T_219_data; // @[RF.scala 32:36]
  wire [63:0] _T_223 = _T_31__T_222_data; // @[RF.scala 32:36]
  wire [63:0] _T_226 = _T_31__T_225_data; // @[RF.scala 32:36]
  wire [63:0] _T_229 = _T_31__T_228_data; // @[RF.scala 32:36]
  wire [63:0] _T_232 = _T_31__T_231_data; // @[RF.scala 32:36]
  wire [63:0] _T_235 = _T_31__T_234_data; // @[RF.scala 32:36]
  wire [63:0] _T_238 = _T_31__T_237_data; // @[RF.scala 32:36]
  wire [63:0] _T_241 = _T_31__T_240_data; // @[RF.scala 32:36]
  wire [63:0] _T_244 = _T_31__T_243_data; // @[RF.scala 32:36]
  wire [63:0] _T_247 = _T_31__T_246_data; // @[RF.scala 32:36]
  wire [63:0] _T_250 = _T_31__T_249_data; // @[RF.scala 32:36]
  wire [63:0] _T_253 = _T_31__T_252_data; // @[RF.scala 32:36]
  wire [63:0] _T_256 = _T_31__T_255_data; // @[RF.scala 32:36]
  wire [63:0] _T_259 = _T_31__T_258_data; // @[RF.scala 32:36]
  wire [63:0] _T_262 = _T_31__T_261_data; // @[RF.scala 32:36]
  wire [63:0] _T_265 = _T_31__T_264_data; // @[RF.scala 32:36]
  wire [63:0] _T_268 = _T_31__T_267_data; // @[RF.scala 32:36]
  wire [63:0] _T_271 = _T_31__T_270_data; // @[RF.scala 32:36]
  wire [63:0] _T_274 = _T_31__T_273_data; // @[RF.scala 32:36]
  wire [63:0] _T_277 = _T_31__T_276_data; // @[RF.scala 32:36]
  wire [63:0] _T_280 = _T_31__T_279_data; // @[RF.scala 32:36]
  wire [63:0] _T_283 = _T_31__T_282_data; // @[RF.scala 32:36]
  wire [63:0] _T_284_0 = 64'h0; // @[ISU.scala 144:34 ISU.scala 144:34]
  wire [63:0] _T_284_1 = _T_193; // @[ISU.scala 144:34 ISU.scala 144:34]
  wire [63:0] _T_284_2 = _T_196; // @[ISU.scala 144:34 ISU.scala 144:34]
  wire [63:0] _T_284_3 = _T_199; // @[ISU.scala 144:34 ISU.scala 144:34]
  wire [63:0] _T_284_4 = _T_202; // @[ISU.scala 144:34 ISU.scala 144:34]
  wire [63:0] _T_284_5 = _T_205; // @[ISU.scala 144:34 ISU.scala 144:34]
  wire [63:0] _T_284_6 = _T_208; // @[ISU.scala 144:34 ISU.scala 144:34]
  wire [63:0] _T_284_7 = _T_211; // @[ISU.scala 144:34 ISU.scala 144:34]
  wire [63:0] _T_284_8 = _T_214; // @[ISU.scala 144:34 ISU.scala 144:34]
  wire [63:0] _T_284_9 = _T_217; // @[ISU.scala 144:34 ISU.scala 144:34]
  wire [63:0] _T_284_10 = _T_220; // @[ISU.scala 144:34 ISU.scala 144:34]
  wire [63:0] _T_284_11 = _T_223; // @[ISU.scala 144:34 ISU.scala 144:34]
  wire [63:0] _T_284_12 = _T_226; // @[ISU.scala 144:34 ISU.scala 144:34]
  wire [63:0] _T_284_13 = _T_229; // @[ISU.scala 144:34 ISU.scala 144:34]
  wire [63:0] _T_284_14 = _T_232; // @[ISU.scala 144:34 ISU.scala 144:34]
  wire [63:0] _T_284_15 = _T_235; // @[ISU.scala 144:34 ISU.scala 144:34]
  wire [63:0] _T_284_16 = _T_238; // @[ISU.scala 144:34 ISU.scala 144:34]
  wire [63:0] _T_284_17 = _T_241; // @[ISU.scala 144:34 ISU.scala 144:34]
  wire [63:0] _T_284_18 = _T_244; // @[ISU.scala 144:34 ISU.scala 144:34]
  wire [63:0] _T_284_19 = _T_247; // @[ISU.scala 144:34 ISU.scala 144:34]
  wire [63:0] _T_284_20 = _T_250; // @[ISU.scala 144:34 ISU.scala 144:34]
  wire [63:0] _T_284_21 = _T_253; // @[ISU.scala 144:34 ISU.scala 144:34]
  wire [63:0] _T_284_22 = _T_256; // @[ISU.scala 144:34 ISU.scala 144:34]
  wire [63:0] _T_284_23 = _T_259; // @[ISU.scala 144:34 ISU.scala 144:34]
  wire [63:0] _T_284_24 = _T_262; // @[ISU.scala 144:34 ISU.scala 144:34]
  wire [63:0] _T_284_25 = _T_265; // @[ISU.scala 144:34 ISU.scala 144:34]
  wire [63:0] _T_284_26 = _T_268; // @[ISU.scala 144:34 ISU.scala 144:34]
  wire [63:0] _T_284_27 = _T_271; // @[ISU.scala 144:34 ISU.scala 144:34]
  wire [63:0] _T_284_28 = _T_274; // @[ISU.scala 144:34 ISU.scala 144:34]
  wire [63:0] _T_284_29 = _T_277; // @[ISU.scala 144:34 ISU.scala 144:34]
  wire [63:0] _T_284_30 = _T_280; // @[ISU.scala 144:34 ISU.scala 144:34]
  wire [63:0] _T_284_31 = _T_283; // @[ISU.scala 144:34 ISU.scala 144:34]
  assign _T_31__T_84_addr = io_in_0_bits_ctrl_rfSrc1;
  assign _T_31__T_84_data = _T_31[_T_31__T_84_addr]; // @[RF.scala 31:15]
  assign _T_31__T_103_addr = io_in_0_bits_ctrl_rfSrc2;
  assign _T_31__T_103_data = _T_31[_T_31__T_103_addr]; // @[RF.scala 31:15]
  assign _T_31__T_189_addr = 5'h0;
  assign _T_31__T_189_data = _T_31[_T_31__T_189_addr]; // @[RF.scala 31:15]
  assign _T_31__T_192_addr = 5'h1;
  assign _T_31__T_192_data = _T_31[_T_31__T_192_addr]; // @[RF.scala 31:15]
  assign _T_31__T_195_addr = 5'h2;
  assign _T_31__T_195_data = _T_31[_T_31__T_195_addr]; // @[RF.scala 31:15]
  assign _T_31__T_198_addr = 5'h3;
  assign _T_31__T_198_data = _T_31[_T_31__T_198_addr]; // @[RF.scala 31:15]
  assign _T_31__T_201_addr = 5'h4;
  assign _T_31__T_201_data = _T_31[_T_31__T_201_addr]; // @[RF.scala 31:15]
  assign _T_31__T_204_addr = 5'h5;
  assign _T_31__T_204_data = _T_31[_T_31__T_204_addr]; // @[RF.scala 31:15]
  assign _T_31__T_207_addr = 5'h6;
  assign _T_31__T_207_data = _T_31[_T_31__T_207_addr]; // @[RF.scala 31:15]
  assign _T_31__T_210_addr = 5'h7;
  assign _T_31__T_210_data = _T_31[_T_31__T_210_addr]; // @[RF.scala 31:15]
  assign _T_31__T_213_addr = 5'h8;
  assign _T_31__T_213_data = _T_31[_T_31__T_213_addr]; // @[RF.scala 31:15]
  assign _T_31__T_216_addr = 5'h9;
  assign _T_31__T_216_data = _T_31[_T_31__T_216_addr]; // @[RF.scala 31:15]
  assign _T_31__T_219_addr = 5'ha;
  assign _T_31__T_219_data = _T_31[_T_31__T_219_addr]; // @[RF.scala 31:15]
  assign _T_31__T_222_addr = 5'hb;
  assign _T_31__T_222_data = _T_31[_T_31__T_222_addr]; // @[RF.scala 31:15]
  assign _T_31__T_225_addr = 5'hc;
  assign _T_31__T_225_data = _T_31[_T_31__T_225_addr]; // @[RF.scala 31:15]
  assign _T_31__T_228_addr = 5'hd;
  assign _T_31__T_228_data = _T_31[_T_31__T_228_addr]; // @[RF.scala 31:15]
  assign _T_31__T_231_addr = 5'he;
  assign _T_31__T_231_data = _T_31[_T_31__T_231_addr]; // @[RF.scala 31:15]
  assign _T_31__T_234_addr = 5'hf;
  assign _T_31__T_234_data = _T_31[_T_31__T_234_addr]; // @[RF.scala 31:15]
  assign _T_31__T_237_addr = 5'h10;
  assign _T_31__T_237_data = _T_31[_T_31__T_237_addr]; // @[RF.scala 31:15]
  assign _T_31__T_240_addr = 5'h11;
  assign _T_31__T_240_data = _T_31[_T_31__T_240_addr]; // @[RF.scala 31:15]
  assign _T_31__T_243_addr = 5'h12;
  assign _T_31__T_243_data = _T_31[_T_31__T_243_addr]; // @[RF.scala 31:15]
  assign _T_31__T_246_addr = 5'h13;
  assign _T_31__T_246_data = _T_31[_T_31__T_246_addr]; // @[RF.scala 31:15]
  assign _T_31__T_249_addr = 5'h14;
  assign _T_31__T_249_data = _T_31[_T_31__T_249_addr]; // @[RF.scala 31:15]
  assign _T_31__T_252_addr = 5'h15;
  assign _T_31__T_252_data = _T_31[_T_31__T_252_addr]; // @[RF.scala 31:15]
  assign _T_31__T_255_addr = 5'h16;
  assign _T_31__T_255_data = _T_31[_T_31__T_255_addr]; // @[RF.scala 31:15]
  assign _T_31__T_258_addr = 5'h17;
  assign _T_31__T_258_data = _T_31[_T_31__T_258_addr]; // @[RF.scala 31:15]
  assign _T_31__T_261_addr = 5'h18;
  assign _T_31__T_261_data = _T_31[_T_31__T_261_addr]; // @[RF.scala 31:15]
  assign _T_31__T_264_addr = 5'h19;
  assign _T_31__T_264_data = _T_31[_T_31__T_264_addr]; // @[RF.scala 31:15]
  assign _T_31__T_267_addr = 5'h1a;
  assign _T_31__T_267_data = _T_31[_T_31__T_267_addr]; // @[RF.scala 31:15]
  assign _T_31__T_270_addr = 5'h1b;
  assign _T_31__T_270_data = _T_31[_T_31__T_270_addr]; // @[RF.scala 31:15]
  assign _T_31__T_273_addr = 5'h1c;
  assign _T_31__T_273_data = _T_31[_T_31__T_273_addr]; // @[RF.scala 31:15]
  assign _T_31__T_276_addr = 5'h1d;
  assign _T_31__T_276_data = _T_31[_T_31__T_276_addr]; // @[RF.scala 31:15]
  assign _T_31__T_279_addr = 5'h1e;
  assign _T_31__T_279_data = _T_31[_T_31__T_279_addr]; // @[RF.scala 31:15]
  assign _T_31__T_282_addr = 5'h1f;
  assign _T_31__T_282_data = _T_31[_T_31__T_282_addr]; // @[RF.scala 31:15]
  assign _T_31__T_113_data = io_wb_rfData;
  assign _T_31__T_113_addr = io_wb_rfDest;
  assign _T_31__T_113_mask = 1'h1;
  assign _T_31__T_113_en = io_wb_rfWen;
  assign _T_32__T_46_addr = 3'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_32__T_46_data = _T_32[_T_32__T_46_addr]; // @[RF.scala 50:16]
  `else
  assign _T_32__T_46_data = _T_32__T_46_addr >= 3'h6 ? _RAND_2[63:0] : _T_32[_T_32__T_46_addr]; // @[RF.scala 50:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_32__T_51_addr = 3'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_32__T_51_data = _T_32[_T_32__T_51_addr]; // @[RF.scala 50:16]
  `else
  assign _T_32__T_51_data = _T_32__T_51_addr >= 3'h6 ? _RAND_3[63:0] : _T_32[_T_32__T_51_addr]; // @[RF.scala 50:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_32__T_56_addr = 3'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_32__T_56_data = _T_32[_T_32__T_56_addr]; // @[RF.scala 50:16]
  `else
  assign _T_32__T_56_data = _T_32__T_56_addr >= 3'h6 ? _RAND_4[63:0] : _T_32[_T_32__T_56_addr]; // @[RF.scala 50:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_32__T_61_addr = 3'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_32__T_61_data = _T_32[_T_32__T_61_addr]; // @[RF.scala 50:16]
  `else
  assign _T_32__T_61_data = _T_32__T_61_addr >= 3'h6 ? _RAND_5[63:0] : _T_32[_T_32__T_61_addr]; // @[RF.scala 50:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_32__T_66_addr = 3'h5;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_32__T_66_data = _T_32[_T_32__T_66_addr]; // @[RF.scala 50:16]
  `else
  assign _T_32__T_66_data = _T_32__T_66_addr >= 3'h6 ? _RAND_6[63:0] : _T_32[_T_32__T_66_addr]; // @[RF.scala 50:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_32__T_118_addr = 3'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_32__T_118_data = _T_32[_T_32__T_118_addr]; // @[RF.scala 50:16]
  `else
  assign _T_32__T_118_data = _T_32__T_118_addr >= 3'h6 ? _RAND_7[63:0] : _T_32[_T_32__T_118_addr]; // @[RF.scala 50:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_32__T_121_addr = 3'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_32__T_121_data = _T_32[_T_32__T_121_addr]; // @[RF.scala 50:16]
  `else
  assign _T_32__T_121_data = _T_32__T_121_addr >= 3'h6 ? _RAND_8[63:0] : _T_32[_T_32__T_121_addr]; // @[RF.scala 50:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_32__T_124_addr = 3'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_32__T_124_data = _T_32[_T_32__T_124_addr]; // @[RF.scala 50:16]
  `else
  assign _T_32__T_124_data = _T_32__T_124_addr >= 3'h6 ? _RAND_9[63:0] : _T_32[_T_32__T_124_addr]; // @[RF.scala 50:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_32__T_127_addr = 3'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_32__T_127_data = _T_32[_T_32__T_127_addr]; // @[RF.scala 50:16]
  `else
  assign _T_32__T_127_data = _T_32__T_127_addr >= 3'h6 ? _RAND_10[63:0] : _T_32[_T_32__T_127_addr]; // @[RF.scala 50:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_32__T_130_addr = 3'h5;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_32__T_130_data = _T_32[_T_32__T_130_addr]; // @[RF.scala 50:16]
  `else
  assign _T_32__T_130_data = _T_32__T_130_addr >= 3'h6 ? _RAND_11[63:0] : _T_32[_T_32__T_130_addr]; // @[RF.scala 50:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_32__T_69_data = io_wb_srfData;
  assign _T_32__T_69_addr = io_wb_srfDest;
  assign _T_32__T_69_mask = 1'h1;
  assign _T_32__T_69_en = io_wb_srfWen;
  assign io_in_0_ready = _T_169 | _T_155; // @[ISU.scala 133:18]
  assign io_out_valid = _T_29 & src2Ready; // @[ISU.scala 59:16]
  assign io_out_bits_cf_instr = io_in_0_bits_cf_instr; // @[ISU.scala 98:18]
  assign io_out_bits_cf_pc = io_in_0_bits_cf_pc; // @[ISU.scala 98:18]
  assign io_out_bits_cf_pnpc = io_in_0_bits_cf_pnpc; // @[ISU.scala 98:18]
  assign io_out_bits_cf_exceptionVec_1 = io_in_0_bits_cf_exceptionVec_1; // @[ISU.scala 98:18]
  assign io_out_bits_cf_exceptionVec_2 = io_in_0_bits_cf_exceptionVec_2; // @[ISU.scala 98:18]
  assign io_out_bits_cf_exceptionVec_12 = io_in_0_bits_cf_exceptionVec_12; // @[ISU.scala 98:18]
  assign io_out_bits_cf_intrVec_0 = io_in_0_bits_cf_intrVec_0; // @[ISU.scala 98:18]
  assign io_out_bits_cf_intrVec_1 = io_in_0_bits_cf_intrVec_1; // @[ISU.scala 98:18]
  assign io_out_bits_cf_intrVec_2 = io_in_0_bits_cf_intrVec_2; // @[ISU.scala 98:18]
  assign io_out_bits_cf_intrVec_3 = io_in_0_bits_cf_intrVec_3; // @[ISU.scala 98:18]
  assign io_out_bits_cf_intrVec_4 = io_in_0_bits_cf_intrVec_4; // @[ISU.scala 98:18]
  assign io_out_bits_cf_intrVec_5 = io_in_0_bits_cf_intrVec_5; // @[ISU.scala 98:18]
  assign io_out_bits_cf_intrVec_6 = io_in_0_bits_cf_intrVec_6; // @[ISU.scala 98:18]
  assign io_out_bits_cf_intrVec_7 = io_in_0_bits_cf_intrVec_7; // @[ISU.scala 98:18]
  assign io_out_bits_cf_intrVec_8 = io_in_0_bits_cf_intrVec_8; // @[ISU.scala 98:18]
  assign io_out_bits_cf_intrVec_9 = io_in_0_bits_cf_intrVec_9; // @[ISU.scala 98:18]
  assign io_out_bits_cf_intrVec_10 = io_in_0_bits_cf_intrVec_10; // @[ISU.scala 98:18]
  assign io_out_bits_cf_intrVec_11 = io_in_0_bits_cf_intrVec_11; // @[ISU.scala 98:18]
  assign io_out_bits_cf_brIdx = io_in_0_bits_cf_brIdx; // @[ISU.scala 98:18]
  assign io_out_bits_cf_crossPageIPFFix = io_in_0_bits_cf_crossPageIPFFix; // @[ISU.scala 98:18]
  assign io_out_bits_ctrl_fuType = io_in_0_bits_ctrl_fuType; // @[ISU.scala 99:20]
  assign io_out_bits_ctrl_fuOpType = io_in_0_bits_ctrl_fuOpType; // @[ISU.scala 99:20]
  assign io_out_bits_ctrl_rfWen = io_in_0_bits_ctrl_rfWen; // @[ISU.scala 99:20]
  assign io_out_bits_ctrl_rfDest = io_in_0_bits_ctrl_rfDest; // @[ISU.scala 99:20]
  assign io_out_bits_ctrl_isNutCoreTrap = io_in_0_bits_ctrl_isNutCoreTrap; // @[ISU.scala 99:20]
  assign io_out_bits_data_src1 = _T_91 | _T_89; // @[ISU.scala 84:25]
  assign io_out_bits_data_src2 = _T_110 | _T_108; // @[ISU.scala 90:25]
  assign io_out_bits_data_imm = io_in_0_bits_data_imm; // @[ISU.scala 96:25]
  assign io_out_bits_data_srf_0 = _T_44 ? io_forward_wb_srfData : _T_67; // @[ISU.scala 79:37]
  assign io_out_bits_data_srf_1 = _T_44 ? io_forward_wb_srfData : _T_47; // @[ISU.scala 71:37 ISU.scala 79:37]
  assign io_out_bits_data_srf_2 = _T_44 ? io_forward_wb_srfData : _T_52; // @[ISU.scala 73:38 ISU.scala 79:37]
  assign io_out_bits_data_srf_3 = _T_44 ? io_forward_wb_srfData : _T_57; // @[ISU.scala 75:37 ISU.scala 79:37]
  assign _T_183_0 = _T_183;
  assign _T_284_0_0 = _T_190;
  assign _T_284_0_1 = _T_284_1;
  assign _T_284_0_2 = _T_284_2;
  assign _T_284_0_3 = _T_284_3;
  assign _T_284_0_4 = _T_284_4;
  assign _T_284_0_5 = _T_284_5;
  assign _T_284_0_6 = _T_284_6;
  assign _T_284_0_7 = _T_284_7;
  assign _T_284_0_8 = _T_284_8;
  assign _T_284_0_9 = _T_284_9;
  assign _T_284_0_10 = _T_284_10;
  assign _T_284_0_11 = _T_284_11;
  assign _T_284_0_12 = _T_284_12;
  assign _T_284_0_13 = _T_284_13;
  assign _T_284_0_14 = _T_284_14;
  assign _T_284_0_15 = _T_284_15;
  assign _T_284_0_16 = _T_284_16;
  assign _T_284_0_17 = _T_284_17;
  assign _T_284_0_18 = _T_284_18;
  assign _T_284_0_19 = _T_284_19;
  assign _T_284_0_20 = _T_284_20;
  assign _T_284_0_21 = _T_284_21;
  assign _T_284_0_22 = _T_284_22;
  assign _T_284_0_23 = _T_284_23;
  assign _T_284_0_24 = _T_284_24;
  assign _T_284_0_25 = _T_284_25;
  assign _T_284_0_26 = _T_284_26;
  assign _T_284_0_27 = _T_284_27;
  assign _T_284_0_28 = _T_284_28;
  assign _T_284_0_29 = _T_284_29;
  assign _T_284_0_30 = _T_284_30;
  assign _T_284_0_31 = _T_284_31;
  assign _T_186_0 = _T_186;
  assign _T_187_0 = _T_155;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_2 = {2{`RANDOM}};
  _RAND_3 = {2{`RANDOM}};
  _RAND_4 = {2{`RANDOM}};
  _RAND_5 = {2{`RANDOM}};
  _RAND_6 = {2{`RANDOM}};
  _RAND_7 = {2{`RANDOM}};
  _RAND_8 = {2{`RANDOM}};
  _RAND_9 = {2{`RANDOM}};
  _RAND_10 = {2{`RANDOM}};
  _RAND_11 = {2{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    _T_31[initvar] = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  for (initvar = 0; initvar < 6; initvar = initvar+1)
    _T_32[initvar] = _RAND_1[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_20 = _RAND_12[31:0];
  _RAND_13 = {2{`RANDOM}};
  _T_173 = _RAND_13[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_31__T_113_en & _T_31__T_113_mask) begin
      _T_31[_T_31__T_113_addr] <= _T_31__T_113_data; // @[RF.scala 31:15]
    end
    if(_T_32__T_69_en & _T_32__T_69_mask) begin
      _T_32[_T_32__T_69_addr] <= _T_32__T_69_data; // @[RF.scala 50:16]
    end
    if (reset) begin
      _T_20 <= 32'h0;
    end else if (io_flush) begin
      _T_20 <= 32'h0;
    end else begin
      _T_20 <= _T_168;
    end
    if (reset) begin
      _T_173 <= 64'h0;
    end else begin
      _T_173 <= _T_175;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_177 & _T_120) begin
          $fwrite(32'h80000002,"[%d] ISU: ",_T_173); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_177 & _T_120) begin
          $fwrite(32'h80000002,"issue: pc %x npc %x instr %x src1 %x src2 %x imm %x\n",io_out_bits_cf_pc,io_out_bits_cf_pnpc,io_out_bits_cf_instr,io_out_bits_data_src1,io_out_bits_data_src2,io_out_bits_data_imm); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ALU(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [63:0] io_in_bits_src1,
  input  [63:0] io_in_bits_src2,
  input  [6:0]  io_in_bits_func,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits,
  input  [63:0] io_cfIn_instr,
  input  [38:0] io_cfIn_pc,
  input  [38:0] io_cfIn_pnpc,
  input  [3:0]  io_cfIn_brIdx,
  output [38:0] io_redirect_target,
  output        io_redirect_valid,
  input  [63:0] io_offset,
  output        _T_272_0,
  output        _T_288_0,
  output        _T_308_0,
  output        _T_243_0_valid,
  output [38:0] _T_243_0_pc,
  output        _T_243_0_isMissPredict,
  output [38:0] _T_243_0_actualTarget,
  output        _T_243_0_actualTaken,
  output [6:0]  _T_243_0_fuOpType,
  output [1:0]  _T_243_0_btbType,
  output        _T_243_0_isRVC,
  output        _T_283_0,
  output        _T_249_0,
  output        _T_266_0,
  input         DISPLAY_ENABLE,
  output        _T_250_1,
  output        _T_310_0,
  output        _T_304_0,
  output        _T_277_0,
  output        _T_298_0,
  output        _T_294_0,
  output        _T_261_0,
  output        _T_306_0,
  output        _T_255_0,
  output        _T_302_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire  isAdderSub = ~io_in_bits_func[6]; // @[ALU.scala 86:20]
  wire [63:0] _T_2 = isAdderSub ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_3 = io_in_bits_src2 ^ _T_2; // @[ALU.scala 87:33]
  wire [64:0] _T_4 = io_in_bits_src1 + _T_3; // @[ALU.scala 87:24]
  wire [64:0] _GEN_0 = {{64'd0}, isAdderSub}; // @[ALU.scala 87:60]
  wire [64:0] adderRes = _T_4 + _GEN_0; // @[ALU.scala 87:60]
  wire [63:0] xorRes = io_in_bits_src1 ^ io_in_bits_src2; // @[ALU.scala 88:21]
  wire  sltu = ~adderRes[64]; // @[ALU.scala 89:14]
  wire  slt = xorRes[63] ^ sltu; // @[ALU.scala 90:28]
  wire [63:0] _T_10 = {32'h0,io_in_bits_src1[31:0]}; // @[Cat.scala 29:58]
  wire [31:0] _T_14 = io_in_bits_src1[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_15 = {_T_14,io_in_bits_src1[31:0]}; // @[Cat.scala 29:58]
  wire  _T_16 = 7'h25 == io_in_bits_func; // @[Mux.scala 80:60]
  wire [63:0] _T_17 = _T_16 ? _T_10 : io_in_bits_src1; // @[Mux.scala 80:57]
  wire  _T_18 = 7'h2d == io_in_bits_func; // @[Mux.scala 80:60]
  wire [63:0] shsrc1 = _T_18 ? _T_15 : _T_17; // @[Mux.scala 80:57]
  wire [5:0] shamt = io_in_bits_func[5] ? {{1'd0}, io_in_bits_src2[4:0]} : io_in_bits_src2[5:0]; // @[ALU.scala 96:18]
  wire [126:0] _GEN_1 = {{63'd0}, shsrc1}; // @[ALU.scala 98:33]
  wire [126:0] _T_23 = _GEN_1 << shamt; // @[ALU.scala 98:33]
  wire [63:0] _T_25 = {63'h0,slt}; // @[Cat.scala 29:58]
  wire [63:0] _T_26 = {63'h0,sltu}; // @[Cat.scala 29:58]
  wire [63:0] _T_27 = shsrc1 >> shamt; // @[ALU.scala 102:32]
  wire [63:0] _T_28 = io_in_bits_src1 | io_in_bits_src2; // @[ALU.scala 103:30]
  wire [63:0] _T_29 = io_in_bits_src1 & io_in_bits_src2; // @[ALU.scala 104:30]
  wire [63:0] _T_30 = _T_18 ? _T_15 : _T_17; // @[ALU.scala 105:32]
  wire [63:0] _T_32 = $signed(_T_30) >>> shamt; // @[ALU.scala 105:49]
  wire  _T_33 = 4'h1 == io_in_bits_func[3:0]; // @[Mux.scala 80:60]
  wire [64:0] _T_34 = _T_33 ? {{1'd0}, _T_23[63:0]} : adderRes; // @[Mux.scala 80:57]
  wire  _T_35 = 4'h2 == io_in_bits_func[3:0]; // @[Mux.scala 80:60]
  wire [64:0] _T_36 = _T_35 ? {{1'd0}, _T_25} : _T_34; // @[Mux.scala 80:57]
  wire  _T_37 = 4'h3 == io_in_bits_func[3:0]; // @[Mux.scala 80:60]
  wire [64:0] _T_38 = _T_37 ? {{1'd0}, _T_26} : _T_36; // @[Mux.scala 80:57]
  wire  _T_39 = 4'h4 == io_in_bits_func[3:0]; // @[Mux.scala 80:60]
  wire [64:0] _T_40 = _T_39 ? {{1'd0}, xorRes} : _T_38; // @[Mux.scala 80:57]
  wire  _T_41 = 4'h5 == io_in_bits_func[3:0]; // @[Mux.scala 80:60]
  wire [64:0] _T_42 = _T_41 ? {{1'd0}, _T_27} : _T_40; // @[Mux.scala 80:57]
  wire  _T_43 = 4'h6 == io_in_bits_func[3:0]; // @[Mux.scala 80:60]
  wire [64:0] _T_44 = _T_43 ? {{1'd0}, _T_28} : _T_42; // @[Mux.scala 80:57]
  wire  _T_45 = 4'h7 == io_in_bits_func[3:0]; // @[Mux.scala 80:60]
  wire [64:0] _T_46 = _T_45 ? {{1'd0}, _T_29} : _T_44; // @[Mux.scala 80:57]
  wire  _T_47 = 4'hd == io_in_bits_func[3:0]; // @[Mux.scala 80:60]
  wire [64:0] res = _T_47 ? {{1'd0}, _T_32} : _T_46; // @[Mux.scala 80:57]
  wire [31:0] _T_52 = res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_53 = {_T_52,res[31:0]}; // @[Cat.scala 29:58]
  wire [64:0] aluRes = io_in_bits_func[5] ? {{1'd0}, _T_53} : res; // @[ALU.scala 107:19]
  wire  _T_54 = |xorRes; // @[ALU.scala 110:56]
  wire  _T_55 = ~_T_54; // @[ALU.scala 110:48]
  wire  isBranch = ~io_in_bits_func[3]; // @[ALU.scala 62:30]
  wire  isBru = io_in_bits_func[4]; // @[ALU.scala 61:31]
  wire  _T_58 = 2'h0 == io_in_bits_func[2:1]; // @[LookupTree.scala 24:34]
  wire  _T_59 = 2'h2 == io_in_bits_func[2:1]; // @[LookupTree.scala 24:34]
  wire  _T_60 = 2'h3 == io_in_bits_func[2:1]; // @[LookupTree.scala 24:34]
  wire  _T_61 = _T_58 & _T_55; // @[Mux.scala 27:72]
  wire  _T_62 = _T_59 & slt; // @[Mux.scala 27:72]
  wire  _T_63 = _T_60 & sltu; // @[Mux.scala 27:72]
  wire  _T_64 = _T_61 | _T_62; // @[Mux.scala 27:72]
  wire  _T_65 = _T_64 | _T_63; // @[Mux.scala 27:72]
  wire  taken = _T_65 ^ io_in_bits_func[0]; // @[ALU.scala 117:72]
  wire [63:0] _GEN_2 = {{25'd0}, io_cfIn_pc}; // @[ALU.scala 118:41]
  wire [63:0] _T_69 = _GEN_2 + io_offset; // @[ALU.scala 118:41]
  wire [64:0] _T_70 = isBranch ? {{1'd0}, _T_69} : adderRes; // @[ALU.scala 118:19]
  wire [38:0] target = _T_70[38:0]; // @[ALU.scala 118:63]
  wire  _T_71 = ~taken; // @[ALU.scala 119:26]
  wire  _T_72 = _T_71 & isBranch; // @[ALU.scala 119:33]
  wire  _T_75 = ~io_cfIn_brIdx[0]; // @[ALU.scala 119:64]
  wire  _T_76 = io_redirect_target != io_cfIn_pnpc; // @[ALU.scala 119:105]
  wire  _T_77 = _T_75 | _T_76; // @[ALU.scala 119:82]
  wire  predictWrong = _T_72 ? io_cfIn_brIdx[0] : _T_77; // @[ALU.scala 119:25]
  wire  isRVC = io_cfIn_instr[1:0] != 2'h3; // @[ALU.scala 120:35]
  wire  _T_80 = io_cfIn_instr[1:0] == 2'h3; // @[ALU.scala 121:29]
  wire  _T_81 = _T_80 | isRVC; // @[ALU.scala 121:41]
  wire  _T_82 = ~io_in_valid; // @[ALU.scala 121:53]
  wire  _T_83 = _T_81 | _T_82; // @[ALU.scala 121:50]
  wire  _T_85 = _T_83 | reset; // @[ALU.scala 121:9]
  wire  _T_86 = ~_T_85; // @[ALU.scala 121:9]
  wire  _T_89 = ~isRVC; // @[ALU.scala 122:55]
  wire  _T_90 = _T_80 != _T_89; // @[ALU.scala 122:51]
  wire  _T_91 = io_in_valid & _T_90; // @[ALU.scala 122:15]
  reg [63:0] _T_92; // @[GTimer.scala 24:20]
  wire [63:0] _T_94 = _T_92 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_96 = _T_91 & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  wire  _T_98 = ~reset; // @[Debug.scala 56:24]
  wire [38:0] _T_104 = io_cfIn_pc + 39'h2; // @[ALU.scala 123:71]
  wire [38:0] _T_106 = io_cfIn_pc + 39'h4; // @[ALU.scala 123:89]
  wire [38:0] _T_107 = isRVC ? _T_104 : _T_106; // @[ALU.scala 123:52]
  wire  _T_109 = io_in_valid & isBru; // @[ALU.scala 125:30]
  wire  _T_110 = _T_109 & predictWrong; // @[ALU.scala 125:39]
  wire [24:0] _T_114 = io_cfIn_pc[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_115 = {_T_114,io_cfIn_pc}; // @[Cat.scala 29:58]
  wire [63:0] _T_117 = _T_115 + 64'h4; // @[ALU.scala 131:71]
  wire [63:0] _T_123 = _T_115 + 64'h2; // @[ALU.scala 131:108]
  wire [63:0] _T_124 = _T_89 ? _T_117 : _T_123; // @[ALU.scala 131:32]
  wire [64:0] _T_125 = isBru ? {{1'd0}, _T_124} : aluRes; // @[ALU.scala 131:21]
  reg [63:0] _T_127; // @[GTimer.scala 24:20]
  wire [63:0] _T_129 = _T_127 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_131 = _T_109 & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  reg [63:0] _T_137; // @[GTimer.scala 24:20]
  wire [63:0] _T_139 = _T_137 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_147 = io_in_bits_func == 7'h58; // @[ALU.scala 135:162]
  wire  _T_148 = io_in_bits_func == 7'h5c; // @[ALU.scala 135:188]
  wire  _T_149 = _T_147 | _T_148; // @[ALU.scala 135:180]
  wire  _T_150 = io_in_bits_func == 7'h5a; // @[ALU.scala 135:214]
  wire  _T_151 = io_in_bits_func == 7'h5e; // @[ALU.scala 135:239]
  reg [63:0] _T_152; // @[GTimer.scala 24:20]
  wire [63:0] _T_154 = _T_152 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_161; // @[GTimer.scala 24:20]
  wire [63:0] _T_163 = _T_161 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_178 = 7'h5c == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_179 = 7'h5e == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_180 = 7'h58 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_181 = 7'h5a == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire [1:0] _T_189 = _T_179 ? 2'h3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_191 = _T_181 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _GEN_3 = {{1'd0}, _T_178}; // @[Mux.scala 27:72]
  wire [1:0] _T_198 = _GEN_3 | _T_189; // @[Mux.scala 27:72]
  wire [1:0] _GEN_4 = {{1'd0}, _T_180}; // @[Mux.scala 27:72]
  wire [1:0] _T_199 = _T_198 | _GEN_4; // @[Mux.scala 27:72]
  wire [1:0] _T_200 = _T_199 | _T_191; // @[Mux.scala 27:72]
  reg [63:0] _T_202; // @[GTimer.scala 24:20]
  wire [63:0] _T_204 = _T_202 + 64'h1; // @[GTimer.scala 25:12]
  reg  _T_243_valid; // @[ALU.scala 158:34]
  reg [38:0] _T_243_pc; // @[ALU.scala 158:34]
  reg  _T_243_isMissPredict; // @[ALU.scala 158:34]
  reg [38:0] _T_243_actualTarget; // @[ALU.scala 158:34]
  reg  _T_243_actualTaken; // @[ALU.scala 158:34]
  reg [6:0] _T_243_fuOpType; // @[ALU.scala 158:34]
  reg [1:0] _T_243_btbType; // @[ALU.scala 158:34]
  reg  _T_243_isRVC; // @[ALU.scala 158:34]
  wire  _T_245 = ~predictWrong; // @[ALU.scala 160:35]
  wire  _T_246 = _T_109 & _T_245; // @[ALU.scala 160:32]
  wire  _T_249 = _T_246 & isBranch; // @[ALU.scala 162:33]
  wire  _T_250 = _T_110 & isBranch; // @[ALU.scala 163:33]
  wire  _T_253 = io_cfIn_pc[2:0] == 3'h0; // @[ALU.scala 164:63]
  wire  _T_254 = _T_250 & _T_253; // @[ALU.scala 164:45]
  wire  _T_255 = _T_254 & isRVC; // @[ALU.scala 164:73]
  wire  _T_261 = _T_254 & _T_89; // @[ALU.scala 165:73]
  wire  _T_264 = io_cfIn_pc[2:0] == 3'h2; // @[ALU.scala 166:63]
  wire  _T_265 = _T_250 & _T_264; // @[ALU.scala 166:45]
  wire  _T_266 = _T_265 & isRVC; // @[ALU.scala 166:73]
  wire  _T_272 = _T_265 & _T_89; // @[ALU.scala 167:73]
  wire  _T_275 = io_cfIn_pc[2:0] == 3'h4; // @[ALU.scala 168:63]
  wire  _T_276 = _T_250 & _T_275; // @[ALU.scala 168:45]
  wire  _T_277 = _T_276 & isRVC; // @[ALU.scala 168:73]
  wire  _T_283 = _T_276 & _T_89; // @[ALU.scala 169:73]
  wire  _T_286 = io_cfIn_pc[2:0] == 3'h6; // @[ALU.scala 170:63]
  wire  _T_287 = _T_250 & _T_286; // @[ALU.scala 170:45]
  wire  _T_288 = _T_287 & isRVC; // @[ALU.scala 170:73]
  wire  _T_294 = _T_287 & _T_89; // @[ALU.scala 171:73]
  wire  _T_298 = _T_246 & _T_149; // @[ALU.scala 172:33]
  wire  _T_302 = _T_110 & _T_149; // @[ALU.scala 173:33]
  wire  _T_304 = _T_246 & _T_150; // @[ALU.scala 174:33]
  wire  _T_306 = _T_110 & _T_150; // @[ALU.scala 175:33]
  wire  _T_308 = _T_246 & _T_151; // @[ALU.scala 176:33]
  wire  _T_310 = _T_110 & _T_151; // @[ALU.scala 177:33]
  assign io_out_valid = io_in_valid; // @[ALU.scala 145:16]
  assign io_out_bits = _T_125[63:0]; // @[ALU.scala 131:15]
  assign io_redirect_target = _T_72 ? _T_107 : target; // @[ALU.scala 123:22]
  assign io_redirect_valid = _T_109 & predictWrong; // @[ALU.scala 125:21]
  assign _T_272_0 = _T_272;
  assign _T_288_0 = _T_288;
  assign _T_308_0 = _T_308;
  assign _T_243_0_valid = _T_243_valid;
  assign _T_243_0_pc = _T_243_pc;
  assign _T_243_0_isMissPredict = _T_243_isMissPredict;
  assign _T_243_0_actualTarget = _T_243_actualTarget;
  assign _T_243_0_actualTaken = _T_243_actualTaken;
  assign _T_243_0_fuOpType = _T_243_fuOpType;
  assign _T_243_0_btbType = _T_243_btbType;
  assign _T_243_0_isRVC = _T_243_isRVC;
  assign _T_283_0 = _T_283;
  assign _T_249_0 = _T_249;
  assign _T_266_0 = _T_266;
  assign _T_250_1 = _T_250;
  assign _T_310_0 = _T_310;
  assign _T_304_0 = _T_304;
  assign _T_277_0 = _T_277;
  assign _T_298_0 = _T_298;
  assign _T_294_0 = _T_294;
  assign _T_261_0 = _T_261;
  assign _T_306_0 = _T_306;
  assign _T_255_0 = _T_255;
  assign _T_302_0 = _T_302;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  _T_92 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  _T_127 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  _T_137 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  _T_152 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  _T_161 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  _T_202 = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  _T_243_valid = _RAND_6[0:0];
  _RAND_7 = {2{`RANDOM}};
  _T_243_pc = _RAND_7[38:0];
  _RAND_8 = {1{`RANDOM}};
  _T_243_isMissPredict = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  _T_243_actualTarget = _RAND_9[38:0];
  _RAND_10 = {1{`RANDOM}};
  _T_243_actualTaken = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _T_243_fuOpType = _RAND_11[6:0];
  _RAND_12 = {1{`RANDOM}};
  _T_243_btbType = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  _T_243_isRVC = _RAND_13[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_92 <= 64'h0;
    end else begin
      _T_92 <= _T_94;
    end
    if (reset) begin
      _T_127 <= 64'h0;
    end else begin
      _T_127 <= _T_129;
    end
    if (reset) begin
      _T_137 <= 64'h0;
    end else begin
      _T_137 <= _T_139;
    end
    if (reset) begin
      _T_152 <= 64'h0;
    end else begin
      _T_152 <= _T_154;
    end
    if (reset) begin
      _T_161 <= 64'h0;
    end else begin
      _T_161 <= _T_163;
    end
    if (reset) begin
      _T_202 <= 64'h0;
    end else begin
      _T_202 <= _T_204;
    end
    _T_243_valid <= io_in_valid & isBru;
    _T_243_pc <= io_cfIn_pc;
    if (_T_72) begin
      _T_243_isMissPredict <= io_cfIn_brIdx[0];
    end else begin
      _T_243_isMissPredict <= _T_77;
    end
    _T_243_actualTarget <= _T_70[38:0];
    _T_243_actualTaken <= _T_65 ^ io_in_bits_func[0];
    _T_243_fuOpType <= io_in_bits_func;
    _T_243_btbType <= _T_199 | _T_191;
    _T_243_isRVC <= io_cfIn_instr[1:0] != 2'h3;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_86) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ALU.scala:121 assert(io.cfIn.instr(1,0) === \"b11\".U || isRVC || !valid)\n"); // @[ALU.scala 121:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_86) begin
          $fatal; // @[ALU.scala 121:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_96 & _T_98) begin
          $fwrite(32'h80000002,"[%d] ALU: ",_T_92); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_96 & _T_98) begin
          $fwrite(32'h80000002,"[ERROR] pc %x inst %x rvc %x\n",io_cfIn_pc,io_cfIn_instr,isRVC); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_131 & _T_98) begin
          $fwrite(32'h80000002,"[%d] ALU: ",_T_127); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_131 & _T_98) begin
          $fwrite(32'h80000002,"tgt %x, valid:%d, npc: %x, pdwrong: %x\n",io_redirect_target,io_redirect_valid,io_cfIn_pnpc,predictWrong); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_131 & _T_98) begin
          $fwrite(32'h80000002,"[%d] ALU: ",_T_137); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_131 & _T_98) begin
          $fwrite(32'h80000002,"taken:%d addrRes:%x src1:%x src2:%x func:%x\n",taken,adderRes,io_in_bits_src1,io_in_bits_src2,io_in_bits_func); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_131 & _T_98) begin
          $fwrite(32'h80000002,"[%d] ALU: ",_T_152); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_131 & _T_98) begin
          $fwrite(32'h80000002,"[BPW] pc %x tgt %x, npc: %x, pdwrong: %x type: %x%x%x%x\n",io_cfIn_pc,io_redirect_target,io_cfIn_pnpc,predictWrong,isBranch,_T_149,_T_150,_T_151); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_98) begin
          $fwrite(32'h80000002,"[%d] ALU: ",_T_161); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_98) begin
          $fwrite(32'h80000002,"valid:%d isBru:%d isBranch:%d \n",io_in_valid,isBru,isBranch); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_131 & _T_98) begin
          $fwrite(32'h80000002,"[%d] ALU: ",_T_202); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_131 & _T_98) begin
          $fwrite(32'h80000002," bpuUpdateReq: valid:%d pc:%x isMissPredict:%d actualTarget:%x actualTaken:%x fuOpType:%x btbType:%x isRVC:%d \n",_T_109,io_cfIn_pc,predictWrong,target,taken,io_in_bits_func,_T_200,isRVC); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module LSExecUnit(
  input         clock,
  input         reset,
  input         io__in_valid,
  input  [63:0] io__in_bits_src1,
  input  [6:0]  io__in_bits_func,
  input         io__out_ready,
  output        io__out_valid,
  output [63:0] io__out_bits,
  input  [63:0] io__wdata,
  input         io__dmem_req_ready,
  output        io__dmem_req_valid,
  output [38:0] io__dmem_req_bits_addr,
  output [2:0]  io__dmem_req_bits_size,
  output [3:0]  io__dmem_req_bits_cmd,
  output [7:0]  io__dmem_req_bits_wmask,
  output [63:0] io__dmem_req_bits_wdata,
  output        io__dmem_resp_ready,
  input         io__dmem_resp_valid,
  input  [63:0] io__dmem_resp_bits_rdata,
  output        io__isMMIO,
  output        io__dtlbPF,
  output        io__loadAddrMisaligned,
  output        io__storeAddrMisaligned,
  output        _T_250_0,
  input         DTLBPF,
  input         DISPLAY_ENABLE,
  input         DTLBENABLE,
  input         ISAMO2,
  output [63:0] io_in_bits_src1,
  input         DTLBFINISH,
  output        _T_258_0,
  output        _T_262_0,
  output        io_isMMIO
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] addrLatch; // @[UnpipelinedLSU.scala 333:26]
  wire  _T_1 = io__in_bits_func == 7'h7b; // @[LSU.scala 60:51]
  wire  _T_2 = io__in_bits_func[3] | _T_1; // @[LSU.scala 60:43]
  wire  isStore = io__in_valid & _T_2; // @[UnpipelinedLSU.scala 334:23]
  wire  _T_3 = ~isStore; // @[UnpipelinedLSU.scala 335:21]
  wire  _T_4 = io__in_bits_func != 7'h3; // @[UnpipelinedLSU.scala 335:39]
  wire  partialLoad = _T_3 & _T_4; // @[UnpipelinedLSU.scala 335:30]
  reg [1:0] state; // @[UnpipelinedLSU.scala 338:22]
  wire  _T_5 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_6 = io__dmem_req_ready & io__dmem_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_7 = _T_6 & DTLBENABLE; // @[UnpipelinedLSU.scala 353:29]
  wire  _T_9 = ~DTLBENABLE; // @[UnpipelinedLSU.scala 354:32]
  wire  _T_10 = _T_6 & _T_9; // @[UnpipelinedLSU.scala 354:29]
  wire  _T_11 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = DTLBFINISH & DTLBPF; // @[UnpipelinedLSU.scala 358:24]
  wire  _T_13 = ~DTLBPF; // @[UnpipelinedLSU.scala 359:27]
  wire  _T_14 = DTLBFINISH & _T_13; // @[UnpipelinedLSU.scala 359:24]
  wire  _T_15 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = io__dmem_resp_ready & io__dmem_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_18 = 2'h3 == state; // @[Conditional.scala 37:30]
  reg [63:0] _T_21; // @[GTimer.scala 24:20]
  wire [63:0] _T_23 = _T_21 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_25 = _T_6 & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  wire  _T_27 = ~reset; // @[Debug.scala 56:24]
  reg [63:0] _T_33; // @[GTimer.scala 24:20]
  wire [63:0] _T_35 = _T_33 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_42 = DTLBFINISH & DTLBENABLE; // @[UnpipelinedLSU.scala 367:20]
  reg [63:0] _T_45; // @[GTimer.scala 24:20]
  wire [63:0] _T_47 = _T_45 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_49 = _T_42 & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  wire [63:0] _T_57 = {io__wdata[7:0],io__wdata[7:0],io__wdata[7:0],io__wdata[7:0],io__wdata[7:0],io__wdata[7:0],io__wdata[7:0],io__wdata[7:0]}; // @[Cat.scala 29:58]
  wire [63:0] _T_60 = {io__wdata[15:0],io__wdata[15:0],io__wdata[15:0],io__wdata[15:0]}; // @[Cat.scala 29:58]
  wire [63:0] _T_62 = {io__wdata[31:0],io__wdata[31:0]}; // @[Cat.scala 29:58]
  wire  _T_63 = 2'h0 == io__in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire  _T_64 = 2'h1 == io__in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire  _T_65 = 2'h2 == io__in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire  _T_66 = 2'h3 == io__in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire [63:0] _T_67 = _T_63 ? _T_57 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_68 = _T_64 ? _T_60 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_69 = _T_65 ? _T_62 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_70 = _T_66 ? io__wdata : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_71 = _T_67 | _T_68; // @[Mux.scala 27:72]
  wire [63:0] _T_72 = _T_71 | _T_69; // @[Mux.scala 27:72]
  wire [1:0] _T_79 = _T_64 ? 2'h3 : 2'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_80 = _T_65 ? 4'hf : 4'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_81 = _T_66 ? 8'hff : 8'h0; // @[Mux.scala 27:72]
  wire [1:0] _GEN_13 = {{1'd0}, _T_63}; // @[Mux.scala 27:72]
  wire [1:0] _T_82 = _GEN_13 | _T_79; // @[Mux.scala 27:72]
  wire [3:0] _GEN_14 = {{2'd0}, _T_82}; // @[Mux.scala 27:72]
  wire [3:0] _T_83 = _GEN_14 | _T_80; // @[Mux.scala 27:72]
  wire [7:0] _GEN_15 = {{4'd0}, _T_83}; // @[Mux.scala 27:72]
  wire [7:0] _T_84 = _GEN_15 | _T_81; // @[Mux.scala 27:72]
  wire [14:0] _GEN_16 = {{7'd0}, _T_84}; // @[UnpipelinedLSU.scala 306:8]
  wire [14:0] reqWmask = _GEN_16 << io__in_bits_src1[2:0]; // @[UnpipelinedLSU.scala 306:8]
  wire  _T_88 = state == 2'h0; // @[UnpipelinedLSU.scala 379:37]
  wire  _T_89 = io__in_valid & _T_88; // @[UnpipelinedLSU.scala 379:27]
  wire  _T_90 = ~io__loadAddrMisaligned; // @[UnpipelinedLSU.scala 379:52]
  wire  _T_91 = _T_89 & _T_90; // @[UnpipelinedLSU.scala 379:49]
  wire  _T_92 = ~io__storeAddrMisaligned; // @[UnpipelinedLSU.scala 379:78]
  wire  _T_94 = state != 2'h0; // @[UnpipelinedLSU.scala 382:40]
  wire  _T_95 = DTLBPF & _T_94; // @[UnpipelinedLSU.scala 382:31]
  wire  _T_96 = _T_95 | io__loadAddrMisaligned; // @[UnpipelinedLSU.scala 382:51]
  wire  _T_97 = _T_96 | io__storeAddrMisaligned; // @[UnpipelinedLSU.scala 382:76]
  wire  _T_98 = state == 2'h3; // @[UnpipelinedLSU.scala 382:134]
  wire  _T_100 = state == 2'h2; // @[UnpipelinedLSU.scala 382:180]
  wire  _T_101 = _T_16 & _T_100; // @[UnpipelinedLSU.scala 382:170]
  wire  _T_102 = partialLoad ? _T_98 : _T_101; // @[UnpipelinedLSU.scala 382:114]
  wire  _T_106 = io__out_ready & io__out_valid; // @[Decoupled.scala 40:37]
  reg [63:0] _T_108; // @[GTimer.scala 24:20]
  wire [63:0] _T_110 = _T_108 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_112 = _T_106 & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  reg [63:0] rdataLatch; // @[UnpipelinedLSU.scala 388:27]
  wire  _T_126 = 3'h0 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_127 = 3'h1 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_128 = 3'h2 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_129 = 3'h3 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_130 = 3'h4 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_131 = 3'h5 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_132 = 3'h6 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_133 = 3'h7 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire [63:0] _T_134 = _T_126 ? rdataLatch : 64'h0; // @[Mux.scala 27:72]
  wire [55:0] _T_135 = _T_127 ? rdataLatch[63:8] : 56'h0; // @[Mux.scala 27:72]
  wire [47:0] _T_136 = _T_128 ? rdataLatch[63:16] : 48'h0; // @[Mux.scala 27:72]
  wire [39:0] _T_137 = _T_129 ? rdataLatch[63:24] : 40'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_138 = _T_130 ? rdataLatch[63:32] : 32'h0; // @[Mux.scala 27:72]
  wire [23:0] _T_139 = _T_131 ? rdataLatch[63:40] : 24'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_140 = _T_132 ? rdataLatch[63:48] : 16'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_141 = _T_133 ? rdataLatch[63:56] : 8'h0; // @[Mux.scala 27:72]
  wire [63:0] _GEN_17 = {{8'd0}, _T_135}; // @[Mux.scala 27:72]
  wire [63:0] _T_142 = _T_134 | _GEN_17; // @[Mux.scala 27:72]
  wire [63:0] _GEN_18 = {{16'd0}, _T_136}; // @[Mux.scala 27:72]
  wire [63:0] _T_143 = _T_142 | _GEN_18; // @[Mux.scala 27:72]
  wire [63:0] _GEN_19 = {{24'd0}, _T_137}; // @[Mux.scala 27:72]
  wire [63:0] _T_144 = _T_143 | _GEN_19; // @[Mux.scala 27:72]
  wire [63:0] _GEN_20 = {{32'd0}, _T_138}; // @[Mux.scala 27:72]
  wire [63:0] _T_145 = _T_144 | _GEN_20; // @[Mux.scala 27:72]
  wire [63:0] _GEN_21 = {{40'd0}, _T_139}; // @[Mux.scala 27:72]
  wire [63:0] _T_146 = _T_145 | _GEN_21; // @[Mux.scala 27:72]
  wire [63:0] _GEN_22 = {{48'd0}, _T_140}; // @[Mux.scala 27:72]
  wire [63:0] _T_147 = _T_146 | _GEN_22; // @[Mux.scala 27:72]
  wire [63:0] _GEN_23 = {{56'd0}, _T_141}; // @[Mux.scala 27:72]
  wire [63:0] rdataSel = _T_147 | _GEN_23; // @[Mux.scala 27:72]
  wire [55:0] _T_168 = rdataSel[7] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_169 = {_T_168,rdataSel[7:0]}; // @[Cat.scala 29:58]
  wire [47:0] _T_173 = rdataSel[15] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_174 = {_T_173,rdataSel[15:0]}; // @[Cat.scala 29:58]
  wire [31:0] _T_178 = rdataSel[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_179 = {_T_178,rdataSel[31:0]}; // @[Cat.scala 29:58]
  wire [63:0] _T_181 = {56'h0,rdataSel[7:0]}; // @[Cat.scala 29:58]
  wire [63:0] _T_183 = {48'h0,rdataSel[15:0]}; // @[Cat.scala 29:58]
  wire [63:0] _T_185 = {32'h0,rdataSel[31:0]}; // @[Cat.scala 29:58]
  wire  _T_186 = 7'h0 == io__in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_187 = 7'h1 == io__in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_188 = 7'h2 == io__in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_189 = 7'h4 == io__in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_190 = 7'h5 == io__in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_191 = 7'h6 == io__in_bits_func; // @[LookupTree.scala 24:34]
  wire [63:0] _T_192 = _T_186 ? _T_169 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_193 = _T_187 ? _T_174 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_194 = _T_188 ? _T_179 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_195 = _T_189 ? _T_181 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_196 = _T_190 ? _T_183 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_197 = _T_191 ? _T_185 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_198 = _T_192 | _T_193; // @[Mux.scala 27:72]
  wire [63:0] _T_199 = _T_198 | _T_194; // @[Mux.scala 27:72]
  wire [63:0] _T_200 = _T_199 | _T_195; // @[Mux.scala 27:72]
  wire [63:0] _T_201 = _T_200 | _T_196; // @[Mux.scala 27:72]
  wire [63:0] rdataPartialLoad = _T_201 | _T_197; // @[Mux.scala 27:72]
  wire  _T_205 = ~io__in_bits_src1[0]; // @[UnpipelinedLSU.scala 416:27]
  wire  _T_207 = io__in_bits_src1[1:0] == 2'h0; // @[UnpipelinedLSU.scala 417:29]
  wire  _T_209 = io__in_bits_src1[2:0] == 3'h0; // @[UnpipelinedLSU.scala 418:29]
  wire  _T_215 = _T_64 & _T_205; // @[Mux.scala 27:72]
  wire  _T_216 = _T_65 & _T_207; // @[Mux.scala 27:72]
  wire  _T_217 = _T_66 & _T_209; // @[Mux.scala 27:72]
  wire  _T_218 = _T_63 | _T_215; // @[Mux.scala 27:72]
  wire  _T_219 = _T_218 | _T_216; // @[Mux.scala 27:72]
  wire  addrAligned = _T_219 | _T_217; // @[Mux.scala 27:72]
  wire  _T_224 = io__in_valid & _T_3; // @[UnpipelinedLSU.scala 429:35]
  wire  _T_225 = ~ISAMO2; // @[UnpipelinedLSU.scala 429:50]
  wire  _T_226 = _T_224 & _T_225; // @[UnpipelinedLSU.scala 429:47]
  wire  _T_227 = ~addrAligned; // @[UnpipelinedLSU.scala 429:60]
  wire  _T_229 = isStore | ISAMO2; // @[UnpipelinedLSU.scala 430:47]
  wire  _T_230 = io__in_valid & _T_229; // @[UnpipelinedLSU.scala 430:35]
  wire  _T_233 = io__loadAddrMisaligned | io__storeAddrMisaligned; // @[UnpipelinedLSU.scala 432:31]
  reg [63:0] _T_234; // @[GTimer.scala 24:20]
  wire [63:0] _T_236 = _T_234 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_238 = _T_233 & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  wire  _T_244 = ~io__dmem_req_bits_cmd[0]; // @[SimpleBus.scala 73:18]
  wire  _T_246 = ~io__dmem_req_bits_cmd[3]; // @[SimpleBus.scala 73:29]
  wire  _T_247 = _T_244 & _T_246; // @[SimpleBus.scala 73:26]
  wire  _T_248 = io__dmem_req_valid & _T_247; // @[SimpleBus.scala 104:29]
  wire  _T_250 = _T_248 & _T_6; // @[UnpipelinedLSU.scala 434:39]
  reg  _T_258; // @[StopWatch.scala 24:20]
  wire  _GEN_9 = _T_248 | _T_258; // @[StopWatch.scala 30:20]
  wire  _T_260 = io__dmem_req_valid & io__dmem_req_bits_cmd[0]; // @[SimpleBus.scala 103:29]
  reg  _T_262; // @[StopWatch.scala 24:20]
  wire  _GEN_11 = _T_260 | _T_262; // @[StopWatch.scala 30:20]
  assign io__out_valid = _T_97 | _T_102; // @[UnpipelinedLSU.scala 382:16]
  assign io__out_bits = partialLoad ? rdataPartialLoad : io__dmem_resp_bits_rdata; // @[UnpipelinedLSU.scala 421:15]
  assign io__dmem_req_valid = _T_91 & _T_92; // @[UnpipelinedLSU.scala 379:18]
  assign io__dmem_req_bits_addr = io__in_bits_src1[38:0]; // @[SimpleBus.scala 64:15]
  assign io__dmem_req_bits_size = {{1'd0}, io__in_bits_func[1:0]}; // @[SimpleBus.scala 66:15]
  assign io__dmem_req_bits_cmd = {{3'd0}, isStore}; // @[SimpleBus.scala 65:14]
  assign io__dmem_req_bits_wmask = reqWmask[7:0]; // @[SimpleBus.scala 68:16]
  assign io__dmem_req_bits_wdata = _T_72 | _T_70; // @[SimpleBus.scala 67:16]
  assign io__dmem_resp_ready = 1'h1; // @[UnpipelinedLSU.scala 380:19]
  assign io__isMMIO = 1'h0;
  assign io__dtlbPF = DTLBPF; // @[UnpipelinedLSU.scala 349:13]
  assign io__loadAddrMisaligned = _T_226 & _T_227; // @[UnpipelinedLSU.scala 429:25]
  assign io__storeAddrMisaligned = _T_230 & _T_227; // @[UnpipelinedLSU.scala 430:26]
  assign _T_250_0 = _T_250;
  assign io_in_bits_src1 = io__in_bits_src1;
  assign _T_258_0 = _T_258;
  assign _T_262_0 = _T_262;
  assign io_isMMIO = io__isMMIO;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  addrLatch = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[1:0];
  _RAND_2 = {2{`RANDOM}};
  _T_21 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  _T_33 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  _T_45 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  _T_108 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  rdataLatch = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  _T_234 = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  _T_258 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _T_262 = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    addrLatch <= io__in_bits_src1;
    if (reset) begin
      state <= 2'h0;
    end else if (_T_5) begin
      if (_T_10) begin
        state <= 2'h2;
      end else if (_T_7) begin
        state <= 2'h1;
      end
    end else if (_T_11) begin
      if (_T_14) begin
        state <= 2'h2;
      end else if (_T_12) begin
        state <= 2'h0;
      end
    end else if (_T_15) begin
      if (_T_16) begin
        if (partialLoad) begin
          state <= 2'h3;
        end else begin
          state <= 2'h0;
        end
      end
    end else if (_T_18) begin
      state <= 2'h0;
    end
    if (reset) begin
      _T_21 <= 64'h0;
    end else begin
      _T_21 <= _T_23;
    end
    if (reset) begin
      _T_33 <= 64'h0;
    end else begin
      _T_33 <= _T_35;
    end
    if (reset) begin
      _T_45 <= 64'h0;
    end else begin
      _T_45 <= _T_47;
    end
    if (reset) begin
      _T_108 <= 64'h0;
    end else begin
      _T_108 <= _T_110;
    end
    rdataLatch <= io__dmem_resp_bits_rdata;
    if (reset) begin
      _T_234 <= 64'h0;
    end else begin
      _T_234 <= _T_236;
    end
    if (reset) begin
      _T_258 <= 1'h0;
    end else if (_T_16) begin
      _T_258 <= 1'h0;
    end else begin
      _T_258 <= _GEN_9;
    end
    if (reset) begin
      _T_262 <= 1'h0;
    end else if (_T_16) begin
      _T_262 <= 1'h0;
    end else begin
      _T_262 <= _GEN_11;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_25 & _T_27) begin
          $fwrite(32'h80000002,"[%d] LSExecUnit: ",_T_21); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_25 & _T_27) begin
          $fwrite(32'h80000002,"[LSU] %x, size %x, wdata_raw %x, isStore %x\n",io__in_bits_src1,io__in_bits_func[1:0],io__wdata,isStore); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_25 & _T_27) begin
          $fwrite(32'h80000002,"[%d] LSExecUnit: ",_T_33); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_25 & _T_27) begin
          $fwrite(32'h80000002,"[LSU] dtlbFinish:%d dtlbEnable:%d dtlbPF:%d state:%d addr:%x dmemReqFire:%d dmemRespFire:%d dmemRdata:%x\n",DTLBFINISH,DTLBENABLE,DTLBPF,state,io__dmem_req_bits_addr,_T_6,_T_16,io__dmem_resp_bits_rdata); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_49 & _T_27) begin
          $fwrite(32'h80000002,"[%d] LSExecUnit: ",_T_45); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_49 & _T_27) begin
          $fwrite(32'h80000002,"[LSU] dtlbFinish:%d dtlbEnable:%d dtlbPF:%d state:%d addr:%x dmemReqFire:%d dmemRespFire:%d dmemRdata:%x\n",DTLBFINISH,DTLBENABLE,DTLBPF,state,io__dmem_req_bits_addr,_T_6,_T_16,io__dmem_resp_bits_rdata); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_112 & _T_27) begin
          $fwrite(32'h80000002,"[%d] LSExecUnit: ",_T_108); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_112 & _T_27) begin
          $fwrite(32'h80000002,"[LSU-EXECUNIT] state %x dresp %x dpf %x lm %x sm %x\n",state,_T_16,DTLBPF,io__loadAddrMisaligned,io__storeAddrMisaligned); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_238 & _T_27) begin
          $fwrite(32'h80000002,"[%d] LSExecUnit: ",_T_234); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_238 & _T_27) begin
          $fwrite(32'h80000002,"misaligned addr detected\n"); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module AtomALU(
  input  [63:0] io_src1,
  input  [63:0] io_src2,
  input  [6:0]  io_func,
  input         io_isWordOp,
  output [63:0] io_result
);
  wire  isAdderSub = ~io_func[6]; // @[LSU.scala 189:20]
  wire [63:0] _T_2 = isAdderSub ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_3 = io_src2 ^ _T_2; // @[LSU.scala 190:33]
  wire [64:0] _T_4 = io_src1 + _T_3; // @[LSU.scala 190:24]
  wire [64:0] _GEN_0 = {{64'd0}, isAdderSub}; // @[LSU.scala 190:60]
  wire [64:0] adderRes = _T_4 + _GEN_0; // @[LSU.scala 190:60]
  wire [63:0] xorRes = io_src1 ^ io_src2; // @[LSU.scala 191:21]
  wire  sltu = ~adderRes[64]; // @[LSU.scala 192:14]
  wire  slt = xorRes[63] ^ sltu; // @[LSU.scala 193:28]
  wire [63:0] _T_9 = io_src1 & io_src2; // @[LSU.scala 199:32]
  wire [63:0] _T_10 = io_src1 | io_src2; // @[LSU.scala 200:32]
  wire [63:0] _T_12 = slt ? io_src1 : io_src2; // @[LSU.scala 201:29]
  wire [63:0] _T_14 = slt ? io_src2 : io_src1; // @[LSU.scala 202:29]
  wire [63:0] _T_16 = sltu ? io_src1 : io_src2; // @[LSU.scala 203:29]
  wire [63:0] _T_18 = sltu ? io_src2 : io_src1; // @[LSU.scala 204:29]
  wire  _T_19 = 6'h22 == io_func[5:0]; // @[Mux.scala 80:60]
  wire [64:0] _T_20 = _T_19 ? {{1'd0}, io_src2} : adderRes; // @[Mux.scala 80:57]
  wire  _T_21 = 6'h24 == io_func[5:0]; // @[Mux.scala 80:60]
  wire [64:0] _T_22 = _T_21 ? {{1'd0}, xorRes} : _T_20; // @[Mux.scala 80:57]
  wire  _T_23 = 6'h25 == io_func[5:0]; // @[Mux.scala 80:60]
  wire [64:0] _T_24 = _T_23 ? {{1'd0}, _T_9} : _T_22; // @[Mux.scala 80:57]
  wire  _T_25 = 6'h26 == io_func[5:0]; // @[Mux.scala 80:60]
  wire [64:0] _T_26 = _T_25 ? {{1'd0}, _T_10} : _T_24; // @[Mux.scala 80:57]
  wire  _T_27 = 6'h37 == io_func[5:0]; // @[Mux.scala 80:60]
  wire [64:0] _T_28 = _T_27 ? {{1'd0}, _T_12} : _T_26; // @[Mux.scala 80:57]
  wire  _T_29 = 6'h30 == io_func[5:0]; // @[Mux.scala 80:60]
  wire [64:0] _T_30 = _T_29 ? {{1'd0}, _T_14} : _T_28; // @[Mux.scala 80:57]
  wire  _T_31 = 6'h31 == io_func[5:0]; // @[Mux.scala 80:60]
  wire [64:0] _T_32 = _T_31 ? {{1'd0}, _T_16} : _T_30; // @[Mux.scala 80:57]
  wire  _T_33 = 6'h32 == io_func[5:0]; // @[Mux.scala 80:60]
  wire [64:0] res = _T_33 ? {{1'd0}, _T_18} : _T_32; // @[Mux.scala 80:57]
  wire [31:0] _T_37 = res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_38 = {_T_37,res[31:0]}; // @[Cat.scala 29:58]
  assign io_result = io_isWordOp ? _T_38 : res[63:0]; // @[LSU.scala 207:13]
endmodule
module UnpipelinedLSU(
  input         clock,
  input         reset,
  output        io__in_ready,
  input         io__in_valid,
  input  [63:0] io__in_bits_src1,
  input  [63:0] io__in_bits_src2,
  input  [6:0]  io__in_bits_func,
  input         io__out_ready,
  output        io__out_valid,
  output [63:0] io__out_bits,
  input  [63:0] io__wdata,
  input  [31:0] io__instr,
  input         io__dmem_req_ready,
  output        io__dmem_req_valid,
  output [38:0] io__dmem_req_bits_addr,
  output [2:0]  io__dmem_req_bits_size,
  output [3:0]  io__dmem_req_bits_cmd,
  output [7:0]  io__dmem_req_bits_wmask,
  output [63:0] io__dmem_req_bits_wdata,
  input         io__dmem_resp_valid,
  input  [63:0] io__dmem_resp_bits_rdata,
  output        io__isMMIO,
  output        io__dtlbPF,
  output        io__loadAddrMisaligned,
  output        io__storeAddrMisaligned,
  output        _T_250,
  output        setLr_0,
  input         DTLBPF,
  input         lsuMMIO_0,
  output        amoReq_0,
  input         DISPLAY_ENABLE,
  input         DTLBENABLE,
  output [63:0] io_in_bits_src1,
  input         DTLBFINISH,
  output        _T_258,
  output [63:0] setLrAddr_0,
  output        _T_262,
  output        io_isMMIO,
  output        setLrVal_0,
  input  [63:0] lr_addr
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  lsExecUnit_clock; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_reset; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__in_valid; // @[UnpipelinedLSU.scala 47:28]
  wire [63:0] lsExecUnit_io__in_bits_src1; // @[UnpipelinedLSU.scala 47:28]
  wire [6:0] lsExecUnit_io__in_bits_func; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__out_ready; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__out_valid; // @[UnpipelinedLSU.scala 47:28]
  wire [63:0] lsExecUnit_io__out_bits; // @[UnpipelinedLSU.scala 47:28]
  wire [63:0] lsExecUnit_io__wdata; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__dmem_req_ready; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__dmem_req_valid; // @[UnpipelinedLSU.scala 47:28]
  wire [38:0] lsExecUnit_io__dmem_req_bits_addr; // @[UnpipelinedLSU.scala 47:28]
  wire [2:0] lsExecUnit_io__dmem_req_bits_size; // @[UnpipelinedLSU.scala 47:28]
  wire [3:0] lsExecUnit_io__dmem_req_bits_cmd; // @[UnpipelinedLSU.scala 47:28]
  wire [7:0] lsExecUnit_io__dmem_req_bits_wmask; // @[UnpipelinedLSU.scala 47:28]
  wire [63:0] lsExecUnit_io__dmem_req_bits_wdata; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__dmem_resp_ready; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__dmem_resp_valid; // @[UnpipelinedLSU.scala 47:28]
  wire [63:0] lsExecUnit_io__dmem_resp_bits_rdata; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__isMMIO; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__dtlbPF; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__loadAddrMisaligned; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__storeAddrMisaligned; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit__T_250_0; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_DTLBPF; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_DISPLAY_ENABLE; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_DTLBENABLE; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_ISAMO2; // @[UnpipelinedLSU.scala 47:28]
  wire [63:0] lsExecUnit_io_in_bits_src1; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_DTLBFINISH; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit__T_258_0; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit__T_262_0; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io_isMMIO; // @[UnpipelinedLSU.scala 47:28]
  wire [63:0] atomALU_io_src1; // @[UnpipelinedLSU.scala 98:25]
  wire [63:0] atomALU_io_src2; // @[UnpipelinedLSU.scala 98:25]
  wire [6:0] atomALU_io_func; // @[UnpipelinedLSU.scala 98:25]
  wire  atomALU_io_isWordOp; // @[UnpipelinedLSU.scala 98:25]
  wire [63:0] atomALU_io_result; // @[UnpipelinedLSU.scala 98:25]
  wire  atomReq = io__in_valid & io__in_bits_func[5]; // @[UnpipelinedLSU.scala 53:26]
  wire  _T_14 = io__in_bits_func == 7'h20; // @[LSU.scala 62:37]
  wire  _T_15 = ~_T_14; // @[LSU.scala 64:49]
  wire  _T_16 = io__in_bits_func[5] & _T_15; // @[LSU.scala 64:46]
  wire  _T_17 = io__in_bits_func == 7'h21; // @[LSU.scala 63:37]
  wire  _T_18 = ~_T_17; // @[LSU.scala 64:64]
  wire  _T_19 = _T_16 & _T_18; // @[LSU.scala 64:61]
  wire  amoReq = io__in_valid & _T_19; // @[UnpipelinedLSU.scala 54:26]
  wire  lrReq = io__in_valid & _T_14; // @[UnpipelinedLSU.scala 55:25]
  wire  scReq = io__in_valid & _T_17; // @[UnpipelinedLSU.scala 56:25]
  wire [2:0] funct3 = io__instr[14:12]; // @[UnpipelinedLSU.scala 64:26]
  wire  _T_23 = io__in_bits_src1 == lr_addr; // @[UnpipelinedLSU.scala 81:28]
  wire  _T_24 = ~_T_23; // @[UnpipelinedLSU.scala 81:21]
  wire  scInvalid = _T_24 & scReq; // @[UnpipelinedLSU.scala 81:40]
  reg [2:0] state; // @[UnpipelinedLSU.scala 95:24]
  reg [63:0] atomMemReg; // @[UnpipelinedLSU.scala 96:25]
  reg [63:0] atomRegReg; // @[UnpipelinedLSU.scala 97:25]
  wire  _T_25 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_28 = ~atomReq; // @[UnpipelinedLSU.scala 141:56]
  wire  _T_29 = io__in_valid & _T_28; // @[UnpipelinedLSU.scala 141:53]
  wire [63:0] _T_31 = io__in_bits_src1 + io__in_bits_src2; // @[UnpipelinedLSU.scala 143:46]
  wire  _T_32 = lsExecUnit_io__out_ready & lsExecUnit_io__out_valid; // @[Decoupled.scala 40:37]
  wire  _T_33 = _T_32 | scInvalid; // @[UnpipelinedLSU.scala 147:66]
  wire  _T_34 = lsExecUnit_io__out_valid | scInvalid; // @[UnpipelinedLSU.scala 148:66]
  wire  _T_36 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_39 = ~amoReq; // @[UnpipelinedLSU.scala 167:28]
  wire  _T_40 = _T_28 | _T_39; // @[UnpipelinedLSU.scala 167:25]
  wire  _T_41 = ~lrReq; // @[UnpipelinedLSU.scala 167:39]
  wire  _T_42 = _T_40 | _T_41; // @[UnpipelinedLSU.scala 167:36]
  wire  _T_43 = ~scReq; // @[UnpipelinedLSU.scala 167:49]
  wire  _T_44 = _T_42 | _T_43; // @[UnpipelinedLSU.scala 167:46]
  wire  _T_46 = _T_44 | reset; // @[UnpipelinedLSU.scala 167:15]
  wire  _T_47 = ~_T_46; // @[UnpipelinedLSU.scala 167:15]
  wire  _T_49 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire [1:0] _T_50 = funct3[0] ? 2'h3 : 2'h2; // @[UnpipelinedLSU.scala 188:42]
  reg [63:0] _T_52; // @[GTimer.scala 24:20]
  wire [63:0] _T_54 = _T_52 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_58 = ~reset; // @[Debug.scala 56:24]
  wire  _T_61 = 3'h6 == state; // @[Conditional.scala 37:30]
  reg [63:0] _T_62; // @[GTimer.scala 24:20]
  wire [63:0] _T_64 = _T_62 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_71 = 3'h7 == state; // @[Conditional.scala 37:30]
  wire [3:0] _T_72 = funct3[0] ? 4'hb : 4'ha; // @[UnpipelinedLSU.scala 219:42]
  reg [63:0] _T_76; // @[GTimer.scala 24:20]
  wire [63:0] _T_78 = _T_76 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_85 = 3'h3 == state; // @[Conditional.scala 37:30]
  reg [63:0] _T_90; // @[GTimer.scala 24:20]
  wire [63:0] _T_92 = _T_90 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_99 = 3'h4 == state; // @[Conditional.scala 37:30]
  reg [63:0] _T_104; // @[GTimer.scala 24:20]
  wire [63:0] _T_106 = _T_104 + 64'h1; // @[GTimer.scala 25:12]
  wire [63:0] _GEN_11 = io__in_bits_src1; // @[Conditional.scala 39:67]
  wire  _GEN_14 = _T_99 & _T_32; // @[Conditional.scala 39:67]
  wire  _GEN_17 = _T_85 | _T_99; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_20 = _T_85 ? {{2'd0}, _T_50} : _T_72; // @[Conditional.scala 39:67]
  wire  _GEN_22 = _T_85 ? _T_32 : _GEN_14; // @[Conditional.scala 39:67]
  wire  _GEN_25 = _T_71 | _GEN_17; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_28 = _T_71 ? _T_72 : _GEN_20; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_29 = _T_71 ? atomMemReg : io__wdata; // @[Conditional.scala 39:67]
  wire  _GEN_30 = _T_71 ? _T_32 : _GEN_22; // @[Conditional.scala 39:67]
  wire  _GEN_33 = _T_61 ? 1'h0 : _GEN_25; // @[Conditional.scala 39:67]
  wire  _GEN_34 = _T_61 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67]
  wire  _GEN_38 = _T_61 ? 1'h0 : _GEN_30; // @[Conditional.scala 39:67]
  wire  _GEN_42 = _T_49 | _GEN_33; // @[Conditional.scala 39:67]
  wire  _GEN_43 = _T_49 | _GEN_34; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_45 = _T_49 ? {{2'd0}, _T_50} : _GEN_28; // @[Conditional.scala 39:67]
  wire  _GEN_47 = _T_49 ? 1'h0 : _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_52 = _T_36 | _GEN_42; // @[Conditional.scala 39:67]
  wire  _GEN_53 = _T_36 | _GEN_43; // @[Conditional.scala 39:67]
  wire [6:0] _GEN_55 = _T_36 ? io__in_bits_func : {{3'd0}, _GEN_45}; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_56 = _T_36 ? io__wdata : _GEN_29; // @[Conditional.scala 39:67]
  wire  _GEN_57 = _T_36 ? _T_32 : _GEN_47; // @[Conditional.scala 39:67]
  wire  _GEN_58 = _T_36 ? lsExecUnit_io__out_valid : _GEN_47; // @[Conditional.scala 39:67]
  wire  _GEN_67 = _T_25 ? _T_33 : _GEN_57; // @[Conditional.scala 40:58]
  wire  _GEN_68 = _T_25 ? _T_34 : _GEN_58; // @[Conditional.scala 40:58]
  wire  _T_113 = DTLBPF | io__loadAddrMisaligned; // @[UnpipelinedLSU.scala 257:17]
  wire  _T_114 = _T_113 | io__storeAddrMisaligned; // @[UnpipelinedLSU.scala 257:42]
  reg [63:0] _T_116; // @[GTimer.scala 24:20]
  wire [63:0] _T_118 = _T_116 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_120 = io__out_valid & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  wire  _T_126 = lrReq | scReq; // @[UnpipelinedLSU.scala 270:38]
  wire  _T_127 = io__out_valid & _T_126; // @[UnpipelinedLSU.scala 270:28]
  wire  _T_128 = state == 3'h7; // @[UnpipelinedLSU.scala 275:52]
  wire [63:0] _T_129 = _T_128 ? atomRegReg : lsExecUnit_io__out_bits; // @[UnpipelinedLSU.scala 275:45]
  reg  mmioReg; // @[UnpipelinedLSU.scala 280:26]
  wire  _T_131 = ~mmioReg; // @[UnpipelinedLSU.scala 281:11]
  wire  setLr = _T_127; // @[UnpipelinedLSU.scala 70:21 UnpipelinedLSU.scala 270:11]
  wire  setLrVal = lrReq; // @[UnpipelinedLSU.scala 71:24 UnpipelinedLSU.scala 271:14]
  wire [63:0] setLrAddr = io__in_bits_src1; // @[UnpipelinedLSU.scala 72:25 UnpipelinedLSU.scala 272:15]
  wire  _GEN_77 = ~_T_25; // @[UnpipelinedLSU.scala 167:15]
  wire  _GEN_78 = _GEN_77 & _T_36; // @[UnpipelinedLSU.scala 167:15]
  wire  _GEN_82 = ~_T_36; // @[Debug.scala 56:24]
  wire  _GEN_83 = _GEN_77 & _GEN_82; // @[Debug.scala 56:24]
  wire  _GEN_84 = _GEN_83 & _T_49; // @[Debug.scala 56:24]
  wire  _GEN_85 = _GEN_84 & _T_32; // @[Debug.scala 56:24]
  wire  _GEN_86 = _GEN_85 & DISPLAY_ENABLE; // @[Debug.scala 56:24]
  wire  _GEN_96 = ~_T_49; // @[Debug.scala 56:24]
  wire  _GEN_97 = _GEN_83 & _GEN_96; // @[Debug.scala 56:24]
  wire  _GEN_98 = _GEN_97 & _T_61; // @[Debug.scala 56:24]
  wire  _GEN_99 = _GEN_98 & DISPLAY_ENABLE; // @[Debug.scala 56:24]
  wire  _GEN_112 = ~_T_61; // @[Debug.scala 56:24]
  wire  _GEN_113 = _GEN_97 & _GEN_112; // @[Debug.scala 56:24]
  wire  _GEN_114 = _GEN_113 & _T_71; // @[Debug.scala 56:24]
  wire  _GEN_115 = _GEN_114 & _T_32; // @[Debug.scala 56:24]
  wire  _GEN_116 = _GEN_115 & DISPLAY_ENABLE; // @[Debug.scala 56:24]
  wire  _GEN_134 = ~_T_71; // @[Debug.scala 56:24]
  wire  _GEN_135 = _GEN_113 & _GEN_134; // @[Debug.scala 56:24]
  wire  _GEN_136 = _GEN_135 & _T_85; // @[Debug.scala 56:24]
  wire  _GEN_137 = _GEN_136 & _T_32; // @[Debug.scala 56:24]
  wire  _GEN_138 = _GEN_137 & DISPLAY_ENABLE; // @[Debug.scala 56:24]
  wire  _GEN_160 = ~_T_85; // @[Debug.scala 56:24]
  wire  _GEN_161 = _GEN_135 & _GEN_160; // @[Debug.scala 56:24]
  wire  _GEN_162 = _GEN_161 & _T_99; // @[Debug.scala 56:24]
  wire  _GEN_163 = _GEN_162 & _T_32; // @[Debug.scala 56:24]
  wire  _GEN_164 = _GEN_163 & DISPLAY_ENABLE; // @[Debug.scala 56:24]
  LSExecUnit lsExecUnit ( // @[UnpipelinedLSU.scala 47:28]
    .clock(lsExecUnit_clock),
    .reset(lsExecUnit_reset),
    .io__in_valid(lsExecUnit_io__in_valid),
    .io__in_bits_src1(lsExecUnit_io__in_bits_src1),
    .io__in_bits_func(lsExecUnit_io__in_bits_func),
    .io__out_ready(lsExecUnit_io__out_ready),
    .io__out_valid(lsExecUnit_io__out_valid),
    .io__out_bits(lsExecUnit_io__out_bits),
    .io__wdata(lsExecUnit_io__wdata),
    .io__dmem_req_ready(lsExecUnit_io__dmem_req_ready),
    .io__dmem_req_valid(lsExecUnit_io__dmem_req_valid),
    .io__dmem_req_bits_addr(lsExecUnit_io__dmem_req_bits_addr),
    .io__dmem_req_bits_size(lsExecUnit_io__dmem_req_bits_size),
    .io__dmem_req_bits_cmd(lsExecUnit_io__dmem_req_bits_cmd),
    .io__dmem_req_bits_wmask(lsExecUnit_io__dmem_req_bits_wmask),
    .io__dmem_req_bits_wdata(lsExecUnit_io__dmem_req_bits_wdata),
    .io__dmem_resp_ready(lsExecUnit_io__dmem_resp_ready),
    .io__dmem_resp_valid(lsExecUnit_io__dmem_resp_valid),
    .io__dmem_resp_bits_rdata(lsExecUnit_io__dmem_resp_bits_rdata),
    .io__isMMIO(lsExecUnit_io__isMMIO),
    .io__dtlbPF(lsExecUnit_io__dtlbPF),
    .io__loadAddrMisaligned(lsExecUnit_io__loadAddrMisaligned),
    .io__storeAddrMisaligned(lsExecUnit_io__storeAddrMisaligned),
    ._T_250_0(lsExecUnit__T_250_0),
    .DTLBPF(lsExecUnit_DTLBPF),
    .DISPLAY_ENABLE(lsExecUnit_DISPLAY_ENABLE),
    .DTLBENABLE(lsExecUnit_DTLBENABLE),
    .ISAMO2(lsExecUnit_ISAMO2),
    .io_in_bits_src1(lsExecUnit_io_in_bits_src1),
    .DTLBFINISH(lsExecUnit_DTLBFINISH),
    ._T_258_0(lsExecUnit__T_258_0),
    ._T_262_0(lsExecUnit__T_262_0),
    .io_isMMIO(lsExecUnit_io_isMMIO)
  );
  AtomALU atomALU ( // @[UnpipelinedLSU.scala 98:25]
    .io_src1(atomALU_io_src1),
    .io_src2(atomALU_io_src2),
    .io_func(atomALU_io_func),
    .io_isWordOp(atomALU_io_isWordOp),
    .io_result(atomALU_io_result)
  );
  assign io__in_ready = _T_114 | _GEN_67; // @[UnpipelinedLSU.scala 126:32 UnpipelinedLSU.scala 136:36 UnpipelinedLSU.scala 147:38 UnpipelinedLSU.scala 165:36 UnpipelinedLSU.scala 190:36 UnpipelinedLSU.scala 207:36 UnpipelinedLSU.scala 221:36 UnpipelinedLSU.scala 235:36 UnpipelinedLSU.scala 249:36 UnpipelinedLSU.scala 260:19]
  assign io__out_valid = _T_114 | _GEN_68; // @[UnpipelinedLSU.scala 125:32 UnpipelinedLSU.scala 137:36 UnpipelinedLSU.scala 148:38 UnpipelinedLSU.scala 166:36 UnpipelinedLSU.scala 191:36 UnpipelinedLSU.scala 208:36 UnpipelinedLSU.scala 222:36 UnpipelinedLSU.scala 236:36 UnpipelinedLSU.scala 250:36 UnpipelinedLSU.scala 259:20]
  assign io__out_bits = scReq ? {{63'd0}, scInvalid} : _T_129; // @[UnpipelinedLSU.scala 275:17]
  assign io__dmem_req_valid = lsExecUnit_io__dmem_req_valid; // @[UnpipelinedLSU.scala 274:13]
  assign io__dmem_req_bits_addr = lsExecUnit_io__dmem_req_bits_addr; // @[UnpipelinedLSU.scala 274:13]
  assign io__dmem_req_bits_size = lsExecUnit_io__dmem_req_bits_size; // @[UnpipelinedLSU.scala 274:13]
  assign io__dmem_req_bits_cmd = lsExecUnit_io__dmem_req_bits_cmd; // @[UnpipelinedLSU.scala 274:13]
  assign io__dmem_req_bits_wmask = lsExecUnit_io__dmem_req_bits_wmask; // @[UnpipelinedLSU.scala 274:13]
  assign io__dmem_req_bits_wdata = lsExecUnit_io__dmem_req_bits_wdata; // @[UnpipelinedLSU.scala 274:13]
  assign io__isMMIO = mmioReg & io__out_valid; // @[UnpipelinedLSU.scala 283:15]
  assign io__dtlbPF = lsExecUnit_io__dtlbPF; // @[UnpipelinedLSU.scala 49:15]
  assign io__loadAddrMisaligned = lsExecUnit_io__loadAddrMisaligned; // @[UnpipelinedLSU.scala 285:27]
  assign io__storeAddrMisaligned = lsExecUnit_io__storeAddrMisaligned; // @[UnpipelinedLSU.scala 286:28]
  assign _T_250 = lsExecUnit__T_250_0;
  assign setLr_0 = setLr;
  assign amoReq_0 = amoReq;
  assign io_in_bits_src1 = lsExecUnit_io_in_bits_src1;
  assign _T_258 = lsExecUnit__T_258_0;
  assign setLrAddr_0 = _GEN_11;
  assign _T_262 = lsExecUnit__T_262_0;
  assign io_isMMIO = lsExecUnit_io_isMMIO;
  assign setLrVal_0 = setLrVal;
  assign lsExecUnit_clock = clock;
  assign lsExecUnit_reset = reset;
  assign lsExecUnit_io__in_valid = _T_25 ? _T_29 : _GEN_52; // @[UnpipelinedLSU.scala 119:32 UnpipelinedLSU.scala 130:36 UnpipelinedLSU.scala 141:38 UnpipelinedLSU.scala 159:36 UnpipelinedLSU.scala 184:36 UnpipelinedLSU.scala 201:36 UnpipelinedLSU.scala 215:36 UnpipelinedLSU.scala 229:36 UnpipelinedLSU.scala 243:36]
  assign lsExecUnit_io__in_bits_src1 = _T_25 ? _T_31 : io__in_bits_src1; // @[UnpipelinedLSU.scala 143:38 UnpipelinedLSU.scala 186:36 UnpipelinedLSU.scala 217:36 UnpipelinedLSU.scala 231:36 UnpipelinedLSU.scala 245:36]
  assign lsExecUnit_io__in_bits_func = _T_25 ? io__in_bits_func : _GEN_55; // @[UnpipelinedLSU.scala 145:38 UnpipelinedLSU.scala 163:36 UnpipelinedLSU.scala 188:36 UnpipelinedLSU.scala 219:36 UnpipelinedLSU.scala 233:36 UnpipelinedLSU.scala 247:36]
  assign lsExecUnit_io__out_ready = _T_25 | _GEN_53; // @[UnpipelinedLSU.scala 142:38 UnpipelinedLSU.scala 160:36 UnpipelinedLSU.scala 185:36 UnpipelinedLSU.scala 202:36 UnpipelinedLSU.scala 216:36 UnpipelinedLSU.scala 230:36 UnpipelinedLSU.scala 244:36]
  assign lsExecUnit_io__wdata = _T_25 ? io__wdata : _GEN_56; // @[UnpipelinedLSU.scala 146:38 UnpipelinedLSU.scala 164:36 UnpipelinedLSU.scala 220:36 UnpipelinedLSU.scala 248:36]
  assign lsExecUnit_io__dmem_req_ready = io__dmem_req_ready; // @[UnpipelinedLSU.scala 274:13]
  assign lsExecUnit_io__dmem_resp_valid = io__dmem_resp_valid; // @[UnpipelinedLSU.scala 274:13]
  assign lsExecUnit_io__dmem_resp_bits_rdata = io__dmem_resp_bits_rdata; // @[UnpipelinedLSU.scala 274:13]
  assign lsExecUnit_DTLBPF = DTLBPF;
  assign lsExecUnit_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign lsExecUnit_DTLBENABLE = DTLBENABLE;
  assign lsExecUnit_ISAMO2 = amoReq;
  assign lsExecUnit_DTLBFINISH = DTLBFINISH;
  assign atomALU_io_src1 = atomMemReg; // @[UnpipelinedLSU.scala 99:21]
  assign atomALU_io_src2 = io__wdata; // @[UnpipelinedLSU.scala 100:21]
  assign atomALU_io_func = io__in_bits_func; // @[UnpipelinedLSU.scala 101:21]
  assign atomALU_io_isWordOp = ~funct3[0]; // @[UnpipelinedLSU.scala 102:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {2{`RANDOM}};
  atomMemReg = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  atomRegReg = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  _T_52 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  _T_62 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  _T_76 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  _T_90 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  _T_104 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  _T_116 = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  mmioReg = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 3'h0;
    end else if (_T_114) begin
      state <= 3'h0;
    end else if (_T_25) begin
      if (scReq) begin
        if (scInvalid) begin
          state <= 3'h0;
        end else begin
          state <= 3'h4;
        end
      end else if (lrReq) begin
        state <= 3'h3;
      end else if (amoReq) begin
        state <= 3'h5;
      end else begin
        state <= 3'h0;
      end
    end else if (_T_36) begin
      if (io__out_valid) begin
        state <= 3'h0;
      end
    end else if (_T_49) begin
      if (_T_32) begin
        state <= 3'h6;
      end
    end else if (_T_61) begin
      state <= 3'h7;
    end else if (_T_71) begin
      if (_T_32) begin
        state <= 3'h0;
      end
    end else if (_T_85) begin
      if (_T_32) begin
        state <= 3'h0;
      end
    end else if (_T_99) begin
      if (_T_32) begin
        state <= 3'h0;
      end
    end
    if (!(_T_25)) begin
      if (!(_T_36)) begin
        if (_T_49) begin
          atomMemReg <= lsExecUnit_io__out_bits;
        end else if (_T_61) begin
          atomMemReg <= atomALU_io_result;
        end
      end
    end
    if (!(_T_25)) begin
      if (!(_T_36)) begin
        if (_T_49) begin
          atomRegReg <= lsExecUnit_io__out_bits;
        end
      end
    end
    if (reset) begin
      _T_52 <= 64'h0;
    end else begin
      _T_52 <= _T_54;
    end
    if (reset) begin
      _T_62 <= 64'h0;
    end else begin
      _T_62 <= _T_64;
    end
    if (reset) begin
      _T_76 <= 64'h0;
    end else begin
      _T_76 <= _T_78;
    end
    if (reset) begin
      _T_90 <= 64'h0;
    end else begin
      _T_90 <= _T_92;
    end
    if (reset) begin
      _T_104 <= 64'h0;
    end else begin
      _T_104 <= _T_106;
    end
    if (reset) begin
      _T_116 <= 64'h0;
    end else begin
      _T_116 <= _T_118;
    end
    if (reset) begin
      mmioReg <= 1'h0;
    end else if (io__out_valid) begin
      mmioReg <= 1'h0;
    end else if (_T_131) begin
      mmioReg <= lsuMMIO_0;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_78 & _T_47) begin
          $fwrite(32'h80000002,"Assertion failed\n    at UnpipelinedLSU.scala:167 assert(!atomReq || !amoReq || !lrReq || !scReq)\n"); // @[UnpipelinedLSU.scala 167:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_78 & _T_47) begin
          $fatal; // @[UnpipelinedLSU.scala 167:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_86 & _T_58) begin
          $fwrite(32'h80000002,"[%d] UnpipelinedLSU: ",_T_52); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_86 & _T_58) begin
          $fwrite(32'h80000002,"[AMO-L] lsExecUnit.io.out.bits %x addr %x src2 %x\n",lsExecUnit_io__out_bits,lsExecUnit_io__in_bits_src1,io__wdata); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_99 & _T_58) begin
          $fwrite(32'h80000002,"[%d] UnpipelinedLSU: ",_T_62); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_99 & _T_58) begin
          $fwrite(32'h80000002,"[AMO-A] src1 %x src2 %x res %x\n",atomMemReg,io__wdata,atomALU_io_result); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_116 & _T_58) begin
          $fwrite(32'h80000002,"[%d] UnpipelinedLSU: ",_T_76); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_116 & _T_58) begin
          $fwrite(32'h80000002,"[AMO-S] atomRegReg %x addr %x\n",atomRegReg,lsExecUnit_io__in_bits_src1); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_138 & _T_58) begin
          $fwrite(32'h80000002,"[%d] UnpipelinedLSU: ",_T_90); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_138 & _T_58) begin
          $fwrite(32'h80000002,"[LR]\n"); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_164 & _T_58) begin
          $fwrite(32'h80000002,"[%d] UnpipelinedLSU: ",_T_104); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_164 & _T_58) begin
          $fwrite(32'h80000002,"[SC] \n"); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_120 & _T_58) begin
          $fwrite(32'h80000002,"[%d] UnpipelinedLSU: ",_T_116); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_120 & _T_58) begin
          $fwrite(32'h80000002,"[LSU-AGU] state %x inv %x inr %x\n",state,io__in_valid,io__in_ready); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Multiplier(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [64:0]  io_in_bits_0,
  input  [64:0]  io_in_bits_1,
  input          io_out_ready,
  output         io_out_valid,
  output [129:0] io_out_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [95:0] _RAND_0;
  reg [95:0] _RAND_1;
  reg [159:0] _RAND_2;
  reg [159:0] _RAND_3;
  reg [159:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  reg [64:0] _T; // @[MDU.scala 56:43]
  reg [64:0] _T_2; // @[MDU.scala 56:43]
  reg [129:0] _T_4; // @[MDU.scala 57:60]
  reg [129:0] _T_5; // @[MDU.scala 57:52]
  reg [129:0] _T_6; // @[MDU.scala 57:44]
  reg  _T_9; // @[MDU.scala 56:43]
  reg  _T_10; // @[MDU.scala 57:60]
  reg  _T_11; // @[MDU.scala 57:52]
  reg  _T_12; // @[MDU.scala 57:44]
  reg  busy; // @[MDU.scala 62:21]
  wire  _T_13 = ~busy; // @[MDU.scala 63:24]
  wire  _T_14 = io_in_valid & _T_13; // @[MDU.scala 63:21]
  wire  _GEN_0 = _T_14 | busy; // @[MDU.scala 63:31]
  assign io_in_ready = ~busy; // @[MDU.scala 65:15]
  assign io_out_valid = _T_12; // @[MDU.scala 60:16]
  assign io_out_bits = _T_6; // @[MDU.scala 59:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {3{`RANDOM}};
  _T = _RAND_0[64:0];
  _RAND_1 = {3{`RANDOM}};
  _T_2 = _RAND_1[64:0];
  _RAND_2 = {5{`RANDOM}};
  _T_4 = _RAND_2[129:0];
  _RAND_3 = {5{`RANDOM}};
  _T_5 = _RAND_3[129:0];
  _RAND_4 = {5{`RANDOM}};
  _T_6 = _RAND_4[129:0];
  _RAND_5 = {1{`RANDOM}};
  _T_9 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _T_10 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_11 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _T_12 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  busy = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T <= io_in_bits_0;
    _T_2 <= io_in_bits_1;
    _T_4 <= $signed(_T) * $signed(_T_2);
    _T_5 <= _T_4;
    _T_6 <= _T_5;
    _T_9 <= io_in_ready & io_in_valid;
    _T_10 <= _T_9;
    _T_11 <= _T_10;
    _T_12 <= _T_11;
    if (reset) begin
      busy <= 1'h0;
    end else if (io_out_valid) begin
      busy <= 1'h0;
    end else begin
      busy <= _GEN_0;
    end
  end
endmodule
module Divider(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [63:0]  io_in_bits_0,
  input  [63:0]  io_in_bits_1,
  input          io_sign,
  output         io_out_valid,
  output [127:0] io_out_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [159:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [95:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[MDU.scala 77:22]
  wire  _T = state == 3'h0; // @[MDU.scala 78:23]
  wire  _T_1 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire  newReq = _T & _T_1; // @[MDU.scala 78:35]
  wire  divBy0 = io_in_bits_1 == 64'h0; // @[MDU.scala 81:18]
  reg [128:0] shiftReg; // @[MDU.scala 83:21]
  wire [64:0] hi = shiftReg[128:64]; // @[MDU.scala 84:20]
  wire [63:0] lo = shiftReg[63:0]; // @[MDU.scala 85:20]
  wire  aSign = io_in_bits_0[63] & io_sign; // @[MDU.scala 72:24]
  wire [63:0] _T_4 = 64'h0 - io_in_bits_0; // @[MDU.scala 73:16]
  wire [63:0] aVal = aSign ? _T_4 : io_in_bits_0; // @[MDU.scala 73:12]
  wire  bSign = io_in_bits_1[63] & io_sign; // @[MDU.scala 72:24]
  wire [63:0] _T_7 = 64'h0 - io_in_bits_1; // @[MDU.scala 73:16]
  reg  aSignReg; // @[Reg.scala 15:16]
  wire  _T_8 = aSign ^ bSign; // @[MDU.scala 90:35]
  wire  _T_9 = ~divBy0; // @[MDU.scala 90:47]
  wire  _T_10 = _T_8 & _T_9; // @[MDU.scala 90:44]
  reg  qSignReg; // @[Reg.scala 15:16]
  reg [63:0] bReg; // @[Reg.scala 15:16]
  wire [64:0] _T_11 = {aVal,1'h0}; // @[Cat.scala 29:58]
  reg [64:0] aValx2Reg; // @[Reg.scala 15:16]
  reg [5:0] value; // @[Counter.scala 29:33]
  wire  _T_12 = state == 3'h1; // @[MDU.scala 97:22]
  wire  _T_15 = |bReg[63:32]; // @[CircuitMath.scala 37:22]
  wire  _T_18 = |bReg[63:48]; // @[CircuitMath.scala 37:22]
  wire  _T_21 = |bReg[63:56]; // @[CircuitMath.scala 37:22]
  wire  _T_24 = |bReg[63:60]; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_28 = bReg[62] ? 2'h2 : {{1'd0}, bReg[61]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_29 = bReg[63] ? 2'h3 : _T_28; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_33 = bReg[58] ? 2'h2 : {{1'd0}, bReg[57]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_34 = bReg[59] ? 2'h3 : _T_33; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_35 = _T_24 ? _T_29 : _T_34; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_36 = {_T_24,_T_35}; // @[Cat.scala 29:58]
  wire  _T_39 = |bReg[55:52]; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_43 = bReg[54] ? 2'h2 : {{1'd0}, bReg[53]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_44 = bReg[55] ? 2'h3 : _T_43; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_48 = bReg[50] ? 2'h2 : {{1'd0}, bReg[49]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_49 = bReg[51] ? 2'h3 : _T_48; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_50 = _T_39 ? _T_44 : _T_49; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_51 = {_T_39,_T_50}; // @[Cat.scala 29:58]
  wire [2:0] _T_52 = _T_21 ? _T_36 : _T_51; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_53 = {_T_21,_T_52}; // @[Cat.scala 29:58]
  wire  _T_56 = |bReg[47:40]; // @[CircuitMath.scala 37:22]
  wire  _T_59 = |bReg[47:44]; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_63 = bReg[46] ? 2'h2 : {{1'd0}, bReg[45]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_64 = bReg[47] ? 2'h3 : _T_63; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_68 = bReg[42] ? 2'h2 : {{1'd0}, bReg[41]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_69 = bReg[43] ? 2'h3 : _T_68; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_70 = _T_59 ? _T_64 : _T_69; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_71 = {_T_59,_T_70}; // @[Cat.scala 29:58]
  wire  _T_74 = |bReg[39:36]; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_78 = bReg[38] ? 2'h2 : {{1'd0}, bReg[37]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_79 = bReg[39] ? 2'h3 : _T_78; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_83 = bReg[34] ? 2'h2 : {{1'd0}, bReg[33]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_84 = bReg[35] ? 2'h3 : _T_83; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_85 = _T_74 ? _T_79 : _T_84; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_86 = {_T_74,_T_85}; // @[Cat.scala 29:58]
  wire [2:0] _T_87 = _T_56 ? _T_71 : _T_86; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_88 = {_T_56,_T_87}; // @[Cat.scala 29:58]
  wire [3:0] _T_89 = _T_18 ? _T_53 : _T_88; // @[CircuitMath.scala 38:21]
  wire [4:0] _T_90 = {_T_18,_T_89}; // @[Cat.scala 29:58]
  wire  _T_93 = |bReg[31:16]; // @[CircuitMath.scala 37:22]
  wire  _T_96 = |bReg[31:24]; // @[CircuitMath.scala 37:22]
  wire  _T_99 = |bReg[31:28]; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_103 = bReg[30] ? 2'h2 : {{1'd0}, bReg[29]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_104 = bReg[31] ? 2'h3 : _T_103; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_108 = bReg[26] ? 2'h2 : {{1'd0}, bReg[25]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_109 = bReg[27] ? 2'h3 : _T_108; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_110 = _T_99 ? _T_104 : _T_109; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_111 = {_T_99,_T_110}; // @[Cat.scala 29:58]
  wire  _T_114 = |bReg[23:20]; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_118 = bReg[22] ? 2'h2 : {{1'd0}, bReg[21]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_119 = bReg[23] ? 2'h3 : _T_118; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_123 = bReg[18] ? 2'h2 : {{1'd0}, bReg[17]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_124 = bReg[19] ? 2'h3 : _T_123; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_125 = _T_114 ? _T_119 : _T_124; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_126 = {_T_114,_T_125}; // @[Cat.scala 29:58]
  wire [2:0] _T_127 = _T_96 ? _T_111 : _T_126; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_128 = {_T_96,_T_127}; // @[Cat.scala 29:58]
  wire  _T_131 = |bReg[15:8]; // @[CircuitMath.scala 37:22]
  wire  _T_134 = |bReg[15:12]; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_138 = bReg[14] ? 2'h2 : {{1'd0}, bReg[13]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_139 = bReg[15] ? 2'h3 : _T_138; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_143 = bReg[10] ? 2'h2 : {{1'd0}, bReg[9]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_144 = bReg[11] ? 2'h3 : _T_143; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_145 = _T_134 ? _T_139 : _T_144; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_146 = {_T_134,_T_145}; // @[Cat.scala 29:58]
  wire  _T_149 = |bReg[7:4]; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_153 = bReg[6] ? 2'h2 : {{1'd0}, bReg[5]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_154 = bReg[7] ? 2'h3 : _T_153; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_158 = bReg[2] ? 2'h2 : {{1'd0}, bReg[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_159 = bReg[3] ? 2'h3 : _T_158; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_160 = _T_149 ? _T_154 : _T_159; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_161 = {_T_149,_T_160}; // @[Cat.scala 29:58]
  wire [2:0] _T_162 = _T_131 ? _T_146 : _T_161; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_163 = {_T_131,_T_162}; // @[Cat.scala 29:58]
  wire [3:0] _T_164 = _T_93 ? _T_128 : _T_163; // @[CircuitMath.scala 38:21]
  wire [4:0] _T_165 = {_T_93,_T_164}; // @[Cat.scala 29:58]
  wire [4:0] _T_166 = _T_15 ? _T_90 : _T_165; // @[CircuitMath.scala 38:21]
  wire [5:0] _T_167 = {_T_15,_T_166}; // @[Cat.scala 29:58]
  wire [6:0] _GEN_18 = {{1'd0}, _T_167}; // @[MDU.scala 105:31]
  wire [6:0] _T_168 = 7'h40 | _GEN_18; // @[MDU.scala 105:31]
  wire  _T_171 = |aValx2Reg[64]; // @[CircuitMath.scala 37:22]
  wire  _T_174 = |aValx2Reg[63:32]; // @[CircuitMath.scala 37:22]
  wire  _T_177 = |aValx2Reg[63:48]; // @[CircuitMath.scala 37:22]
  wire  _T_180 = |aValx2Reg[63:56]; // @[CircuitMath.scala 37:22]
  wire  _T_183 = |aValx2Reg[63:60]; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_187 = aValx2Reg[62] ? 2'h2 : {{1'd0}, aValx2Reg[61]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_188 = aValx2Reg[63] ? 2'h3 : _T_187; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_192 = aValx2Reg[58] ? 2'h2 : {{1'd0}, aValx2Reg[57]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_193 = aValx2Reg[59] ? 2'h3 : _T_192; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_194 = _T_183 ? _T_188 : _T_193; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_195 = {_T_183,_T_194}; // @[Cat.scala 29:58]
  wire  _T_198 = |aValx2Reg[55:52]; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_202 = aValx2Reg[54] ? 2'h2 : {{1'd0}, aValx2Reg[53]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_203 = aValx2Reg[55] ? 2'h3 : _T_202; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_207 = aValx2Reg[50] ? 2'h2 : {{1'd0}, aValx2Reg[49]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_208 = aValx2Reg[51] ? 2'h3 : _T_207; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_209 = _T_198 ? _T_203 : _T_208; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_210 = {_T_198,_T_209}; // @[Cat.scala 29:58]
  wire [2:0] _T_211 = _T_180 ? _T_195 : _T_210; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_212 = {_T_180,_T_211}; // @[Cat.scala 29:58]
  wire  _T_215 = |aValx2Reg[47:40]; // @[CircuitMath.scala 37:22]
  wire  _T_218 = |aValx2Reg[47:44]; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_222 = aValx2Reg[46] ? 2'h2 : {{1'd0}, aValx2Reg[45]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_223 = aValx2Reg[47] ? 2'h3 : _T_222; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_227 = aValx2Reg[42] ? 2'h2 : {{1'd0}, aValx2Reg[41]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_228 = aValx2Reg[43] ? 2'h3 : _T_227; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_229 = _T_218 ? _T_223 : _T_228; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_230 = {_T_218,_T_229}; // @[Cat.scala 29:58]
  wire  _T_233 = |aValx2Reg[39:36]; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_237 = aValx2Reg[38] ? 2'h2 : {{1'd0}, aValx2Reg[37]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_238 = aValx2Reg[39] ? 2'h3 : _T_237; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_242 = aValx2Reg[34] ? 2'h2 : {{1'd0}, aValx2Reg[33]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_243 = aValx2Reg[35] ? 2'h3 : _T_242; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_244 = _T_233 ? _T_238 : _T_243; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_245 = {_T_233,_T_244}; // @[Cat.scala 29:58]
  wire [2:0] _T_246 = _T_215 ? _T_230 : _T_245; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_247 = {_T_215,_T_246}; // @[Cat.scala 29:58]
  wire [3:0] _T_248 = _T_177 ? _T_212 : _T_247; // @[CircuitMath.scala 38:21]
  wire [4:0] _T_249 = {_T_177,_T_248}; // @[Cat.scala 29:58]
  wire  _T_252 = |aValx2Reg[31:16]; // @[CircuitMath.scala 37:22]
  wire  _T_255 = |aValx2Reg[31:24]; // @[CircuitMath.scala 37:22]
  wire  _T_258 = |aValx2Reg[31:28]; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_262 = aValx2Reg[30] ? 2'h2 : {{1'd0}, aValx2Reg[29]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_263 = aValx2Reg[31] ? 2'h3 : _T_262; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_267 = aValx2Reg[26] ? 2'h2 : {{1'd0}, aValx2Reg[25]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_268 = aValx2Reg[27] ? 2'h3 : _T_267; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_269 = _T_258 ? _T_263 : _T_268; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_270 = {_T_258,_T_269}; // @[Cat.scala 29:58]
  wire  _T_273 = |aValx2Reg[23:20]; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_277 = aValx2Reg[22] ? 2'h2 : {{1'd0}, aValx2Reg[21]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_278 = aValx2Reg[23] ? 2'h3 : _T_277; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_282 = aValx2Reg[18] ? 2'h2 : {{1'd0}, aValx2Reg[17]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_283 = aValx2Reg[19] ? 2'h3 : _T_282; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_284 = _T_273 ? _T_278 : _T_283; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_285 = {_T_273,_T_284}; // @[Cat.scala 29:58]
  wire [2:0] _T_286 = _T_255 ? _T_270 : _T_285; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_287 = {_T_255,_T_286}; // @[Cat.scala 29:58]
  wire  _T_290 = |aValx2Reg[15:8]; // @[CircuitMath.scala 37:22]
  wire  _T_293 = |aValx2Reg[15:12]; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_297 = aValx2Reg[14] ? 2'h2 : {{1'd0}, aValx2Reg[13]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_298 = aValx2Reg[15] ? 2'h3 : _T_297; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_302 = aValx2Reg[10] ? 2'h2 : {{1'd0}, aValx2Reg[9]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_303 = aValx2Reg[11] ? 2'h3 : _T_302; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_304 = _T_293 ? _T_298 : _T_303; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_305 = {_T_293,_T_304}; // @[Cat.scala 29:58]
  wire  _T_308 = |aValx2Reg[7:4]; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_312 = aValx2Reg[6] ? 2'h2 : {{1'd0}, aValx2Reg[5]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_313 = aValx2Reg[7] ? 2'h3 : _T_312; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_317 = aValx2Reg[2] ? 2'h2 : {{1'd0}, aValx2Reg[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_318 = aValx2Reg[3] ? 2'h3 : _T_317; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_319 = _T_308 ? _T_313 : _T_318; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_320 = {_T_308,_T_319}; // @[Cat.scala 29:58]
  wire [2:0] _T_321 = _T_290 ? _T_305 : _T_320; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_322 = {_T_290,_T_321}; // @[Cat.scala 29:58]
  wire [3:0] _T_323 = _T_252 ? _T_287 : _T_322; // @[CircuitMath.scala 38:21]
  wire [4:0] _T_324 = {_T_252,_T_323}; // @[Cat.scala 29:58]
  wire [4:0] _T_325 = _T_174 ? _T_249 : _T_324; // @[CircuitMath.scala 38:21]
  wire [5:0] _T_326 = {_T_174,_T_325}; // @[Cat.scala 29:58]
  wire [5:0] _T_327 = _T_171 ? 6'h0 : _T_326; // @[CircuitMath.scala 38:21]
  wire [6:0] _T_328 = {_T_171,_T_327}; // @[Cat.scala 29:58]
  wire [6:0] _T_330 = _T_168 - _T_328; // @[MDU.scala 105:45]
  wire  _T_331 = _T_330 >= 7'h3f; // @[MDU.scala 109:52]
  wire [6:0] _T_332 = _T_331 ? 7'h3f : _T_330; // @[MDU.scala 109:38]
  wire [6:0] _T_333 = divBy0 ? 7'h0 : _T_332; // @[MDU.scala 109:21]
  wire  _T_334 = state == 3'h2; // @[MDU.scala 111:22]
  wire [127:0] _GEN_19 = {{63'd0}, aValx2Reg}; // @[MDU.scala 112:27]
  wire [127:0] _T_335 = _GEN_19 << value; // @[MDU.scala 112:27]
  wire  _T_336 = state == 3'h3; // @[MDU.scala 114:22]
  wire [64:0] _GEN_20 = {{1'd0}, bReg}; // @[MDU.scala 115:28]
  wire  _T_337 = hi >= _GEN_20; // @[MDU.scala 115:28]
  wire [64:0] _T_339 = hi - _GEN_20; // @[MDU.scala 116:36]
  wire [64:0] _T_340 = _T_337 ? _T_339 : hi; // @[MDU.scala 116:24]
  wire [128:0] _T_343 = {_T_340[63:0],lo,_T_337}; // @[Cat.scala 29:58]
  wire  _T_344 = value == 6'h3f; // @[Counter.scala 38:24]
  wire [5:0] _T_346 = value + 6'h1; // @[Counter.scala 39:22]
  wire  _T_348 = state == 3'h4; // @[MDU.scala 119:22]
  wire [5:0] _GEN_7 = _T_336 ? _T_346 : value; // @[MDU.scala 114:37]
  wire [5:0] _GEN_11 = _T_334 ? value : _GEN_7; // @[MDU.scala 111:35]
  wire [6:0] _GEN_12 = _T_12 ? _T_333 : {{1'd0}, _GEN_11}; // @[MDU.scala 97:34]
  wire [6:0] _GEN_16 = newReq ? {{1'd0}, value} : _GEN_12; // @[MDU.scala 95:17]
  wire [63:0] r = hi[64:1]; // @[MDU.scala 123:13]
  wire [63:0] _T_350 = 64'h0 - lo; // @[MDU.scala 124:28]
  wire [63:0] resQ = qSignReg ? _T_350 : lo; // @[MDU.scala 124:17]
  wire [63:0] _T_352 = 64'h0 - r; // @[MDU.scala 125:28]
  wire [63:0] resR = aSignReg ? _T_352 : r; // @[MDU.scala 125:17]
  assign io_in_ready = state == 3'h0; // @[MDU.scala 129:15]
  assign io_out_valid = state == 3'h4; // @[MDU.scala 128:16]
  assign io_out_bits = {resR,resQ}; // @[MDU.scala 126:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {5{`RANDOM}};
  shiftReg = _RAND_1[128:0];
  _RAND_2 = {1{`RANDOM}};
  aSignReg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  qSignReg = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  bReg = _RAND_4[63:0];
  _RAND_5 = {3{`RANDOM}};
  aValx2Reg = _RAND_5[64:0];
  _RAND_6 = {1{`RANDOM}};
  value = _RAND_6[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 3'h0;
    end else if (newReq) begin
      state <= 3'h1;
    end else if (_T_12) begin
      state <= 3'h2;
    end else if (_T_334) begin
      state <= 3'h3;
    end else if (_T_336) begin
      if (_T_344) begin
        state <= 3'h4;
      end
    end else if (_T_348) begin
      state <= 3'h0;
    end
    if (!(newReq)) begin
      if (!(_T_12)) begin
        if (_T_334) begin
          shiftReg <= {{1'd0}, _T_335};
        end else if (_T_336) begin
          shiftReg <= _T_343;
        end
      end
    end
    if (newReq) begin
      aSignReg <= aSign;
    end
    if (newReq) begin
      qSignReg <= _T_10;
    end
    if (newReq) begin
      if (bSign) begin
        bReg <= _T_7;
      end else begin
        bReg <= io_in_bits_1;
      end
    end
    if (newReq) begin
      aValx2Reg <= _T_11;
    end
    if (reset) begin
      value <= 6'h0;
    end else begin
      value <= _GEN_16[5:0];
    end
  end
endmodule
module MDU(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [63:0] io_in_bits_src1,
  input  [63:0] io_in_bits_src2,
  input  [6:0]  io_in_bits_func,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits,
  input         DISPLAY_ENABLE,
  output        _T_87_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  mul_clock; // @[MDU.scala 151:19]
  wire  mul_reset; // @[MDU.scala 151:19]
  wire  mul_io_in_ready; // @[MDU.scala 151:19]
  wire  mul_io_in_valid; // @[MDU.scala 151:19]
  wire [64:0] mul_io_in_bits_0; // @[MDU.scala 151:19]
  wire [64:0] mul_io_in_bits_1; // @[MDU.scala 151:19]
  wire  mul_io_out_ready; // @[MDU.scala 151:19]
  wire  mul_io_out_valid; // @[MDU.scala 151:19]
  wire [129:0] mul_io_out_bits; // @[MDU.scala 151:19]
  wire  div_clock; // @[MDU.scala 152:19]
  wire  div_reset; // @[MDU.scala 152:19]
  wire  div_io_in_ready; // @[MDU.scala 152:19]
  wire  div_io_in_valid; // @[MDU.scala 152:19]
  wire [63:0] div_io_in_bits_0; // @[MDU.scala 152:19]
  wire [63:0] div_io_in_bits_1; // @[MDU.scala 152:19]
  wire  div_io_sign; // @[MDU.scala 152:19]
  wire  div_io_out_valid; // @[MDU.scala 152:19]
  wire [127:0] div_io_out_bits; // @[MDU.scala 152:19]
  wire  isDiv = io_in_bits_func[2]; // @[MDU.scala 41:27]
  wire  _T_2 = ~io_in_bits_func[0]; // @[MDU.scala 42:42]
  wire  isDivSign = isDiv & _T_2; // @[MDU.scala 42:39]
  wire  isW = io_in_bits_func[3]; // @[MDU.scala 43:25]
  wire [64:0] _T_4 = {1'h0,io_in_bits_src1}; // @[Cat.scala 29:58]
  wire [64:0] _T_6 = {io_in_bits_src1[63],io_in_bits_src1}; // @[Cat.scala 29:58]
  wire  _T_10 = 2'h0 == io_in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire  _T_11 = 2'h1 == io_in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire  _T_12 = 2'h2 == io_in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire  _T_13 = 2'h3 == io_in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire [64:0] _T_14 = _T_10 ? _T_4 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_15 = _T_11 ? _T_6 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_16 = _T_12 ? _T_6 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_17 = _T_13 ? _T_4 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_18 = _T_14 | _T_15; // @[Mux.scala 27:72]
  wire [64:0] _T_19 = _T_18 | _T_16; // @[Mux.scala 27:72]
  wire [64:0] _T_23 = {1'h0,io_in_bits_src2}; // @[Cat.scala 29:58]
  wire [64:0] _T_25 = {io_in_bits_src2[63],io_in_bits_src2}; // @[Cat.scala 29:58]
  wire [64:0] _T_32 = _T_10 ? _T_23 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_33 = _T_11 ? _T_25 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_34 = _T_12 ? _T_23 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_35 = _T_13 ? _T_23 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_36 = _T_32 | _T_33; // @[Mux.scala 27:72]
  wire [64:0] _T_37 = _T_36 | _T_34; // @[Mux.scala 27:72]
  wire [31:0] _T_43 = io_in_bits_src1[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_44 = {_T_43,io_in_bits_src1[31:0]}; // @[Cat.scala 29:58]
  wire [63:0] _T_46 = {32'h0,io_in_bits_src1[31:0]}; // @[Cat.scala 29:58]
  wire [63:0] _T_47 = isDivSign ? _T_44 : _T_46; // @[MDU.scala 169:47]
  wire [31:0] _T_52 = io_in_bits_src2[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_53 = {_T_52,io_in_bits_src2[31:0]}; // @[Cat.scala 29:58]
  wire [63:0] _T_55 = {32'h0,io_in_bits_src2[31:0]}; // @[Cat.scala 29:58]
  wire [63:0] _T_56 = isDivSign ? _T_53 : _T_55; // @[MDU.scala 169:47]
  wire  _T_58 = ~isDiv; // @[MDU.scala 173:37]
  wire  _T_62 = io_in_bits_func[1:0] == 2'h0; // @[MDU.scala 176:30]
  wire [63:0] mulRes = _T_62 ? mul_io_out_bits[63:0] : mul_io_out_bits[127:64]; // @[MDU.scala 176:19]
  wire [63:0] divRes = io_in_bits_func[1] ? div_io_out_bits[127:64] : div_io_out_bits[63:0]; // @[MDU.scala 177:19]
  wire [63:0] res = isDiv ? divRes : mulRes; // @[MDU.scala 178:16]
  wire [31:0] _T_71 = res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_72 = {_T_71,res[31:0]}; // @[Cat.scala 29:58]
  wire  _T_74 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  reg  _T_75; // @[MDU.scala 181:50]
  wire  isDivReg = _T_74 ? isDiv : _T_75; // @[MDU.scala 181:21]
  reg [63:0] _T_78; // @[GTimer.scala 24:20]
  wire [63:0] _T_80 = _T_78 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_84 = ~reset; // @[Debug.scala 56:24]
  wire  _T_87 = mul_io_out_ready & mul_io_out_valid; // @[Decoupled.scala 40:37]
  Multiplier mul ( // @[MDU.scala 151:19]
    .clock(mul_clock),
    .reset(mul_reset),
    .io_in_ready(mul_io_in_ready),
    .io_in_valid(mul_io_in_valid),
    .io_in_bits_0(mul_io_in_bits_0),
    .io_in_bits_1(mul_io_in_bits_1),
    .io_out_ready(mul_io_out_ready),
    .io_out_valid(mul_io_out_valid),
    .io_out_bits(mul_io_out_bits)
  );
  Divider div ( // @[MDU.scala 152:19]
    .clock(div_clock),
    .reset(div_reset),
    .io_in_ready(div_io_in_ready),
    .io_in_valid(div_io_in_valid),
    .io_in_bits_0(div_io_in_bits_0),
    .io_in_bits_1(div_io_in_bits_1),
    .io_sign(div_io_sign),
    .io_out_valid(div_io_out_valid),
    .io_out_bits(div_io_out_bits)
  );
  assign io_in_ready = isDiv ? div_io_in_ready : mul_io_in_ready; // @[MDU.scala 182:15]
  assign io_out_valid = isDivReg ? div_io_out_valid : mul_io_out_valid; // @[MDU.scala 183:16]
  assign io_out_bits = isW ? _T_72 : res; // @[MDU.scala 179:15]
  assign _T_87_0 = _T_87;
  assign mul_clock = clock;
  assign mul_reset = reset;
  assign mul_io_in_valid = io_in_valid & _T_58; // @[MDU.scala 173:19]
  assign mul_io_in_bits_0 = _T_19 | _T_17; // @[MDU.scala 166:21]
  assign mul_io_in_bits_1 = _T_37 | _T_35; // @[MDU.scala 167:21]
  assign mul_io_out_ready = 1'h1; // @[MDU.scala 155:17]
  assign div_clock = clock;
  assign div_reset = reset;
  assign div_io_in_valid = io_in_valid & isDiv; // @[MDU.scala 174:19]
  assign div_io_in_bits_0 = isW ? _T_47 : io_in_bits_src1; // @[MDU.scala 170:21]
  assign div_io_in_bits_1 = isW ? _T_56 : io_in_bits_src2; // @[MDU.scala 171:21]
  assign div_io_sign = isDiv & _T_2; // @[MDU.scala 154:12]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_75 = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  _T_78 = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_75 <= io_in_bits_func[2];
    if (reset) begin
      _T_78 <= 64'h0;
    end else begin
      _T_78 <= _T_80;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_84) begin
          $fwrite(32'h80000002,"[%d] MDU: ",_T_78); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_84) begin
          $fwrite(32'h80000002,"[FU-MDU] irv-orv %d %d - %d %d\n",io_in_ready,io_in_valid,1'h1,io_out_valid); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CSR(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [63:0] io_in_bits_src1,
  input  [63:0] io_in_bits_src2,
  input  [6:0]  io_in_bits_func,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits,
  input  [63:0] io_cfIn_instr,
  input  [38:0] io_cfIn_pc,
  input         io_cfIn_exceptionVec_1,
  input         io_cfIn_exceptionVec_2,
  input         io_cfIn_exceptionVec_4,
  input         io_cfIn_exceptionVec_6,
  input         io_cfIn_exceptionVec_12,
  input         io_cfIn_intrVec_0,
  input         io_cfIn_intrVec_1,
  input         io_cfIn_intrVec_2,
  input         io_cfIn_intrVec_3,
  input         io_cfIn_intrVec_4,
  input         io_cfIn_intrVec_5,
  input         io_cfIn_intrVec_6,
  input         io_cfIn_intrVec_7,
  input         io_cfIn_intrVec_8,
  input         io_cfIn_intrVec_9,
  input         io_cfIn_intrVec_10,
  input         io_cfIn_intrVec_11,
  input         io_cfIn_crossPageIPFFix,
  output [38:0] io_redirect_target,
  output        io_redirect_valid,
  input         io_instrValid,
  output [63:0] io_intrNO,
  output [1:0]  io_imemMMU_priviledgeMode,
  output [1:0]  io_dmemMMU_priviledgeMode,
  output        io_dmemMMU_status_sum,
  output        io_dmemMMU_status_mxr,
  input         io_dmemMMU_loadPF,
  input         io_dmemMMU_storePF,
  input  [38:0] io_dmemMMU_addr,
  output        io_wenFix,
  output [63:0] _T_4181_0,
  input         perfCntCondMloadInstr,
  output [63:0] _T_4184_0,
  input         perfCntCondMlsuInstr,
  input         set_lr,
  input         perfCntCondMrawStall,
  input         Custom4,
  input         Custom7,
  output [63:0] _T_4185_0,
  input         MbpRRight,
  output [63:0] perfCnts_2_0,
  output [63:0] satp_0,
  output [1:0]  _T_4178_0,
  input         Custom6,
  input         perfCntCondMinstret,
  input         MbpBRight,
  input         perfCntCondMexuBusy,
  input         perfCntCondMmduInstr,
  input         mtip_0,
  input         Custom3,
  input         DISPLAY_ENABLE,
  input         MbpBWrong,
  input         MbpRWrong,
  input         meip_0,
  input         perfCntCondISUIssue,
  input         nutcoretrap_0,
  input         MbpIRight,
  input         perfCntCondMcsrInstr,
  input         perfCntCondMsnnInstr,
  input         perfCntCondMmulInstr,
  input  [63:0] LSUADDR,
  input         Custom5,
  input         MbpJRight,
  input         perfCntCondMbruInstr,
  output [11:0] intrVec_0,
  input         perfCntCondMaluInstr,
  input         Custom8,
  input         perfCntCondMloadStall,
  input         Custom2,
  input         msip_0,
  input         MbpIWrong,
  input  [63:0] set_lr_addr,
  input         perfCntCondMimemStall,
  input         perfCntCondMstoreStall,
  output [63:0] _T_4183_0,
  output [63:0] _T_4182_0,
  output [63:0] perfCnts_0_0,
  input         perfCntCondMifuFlush,
  output [63:0] _T_4179_0,
  input         perfCntCondMmmioInstr,
  input         perfCntCondMultiCommit,
  input         Custom1,
  input         MbpJWrong,
  input         set_lr_val,
  output [63:0] lrAddr_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [63:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [63:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [63:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [63:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [63:0] _RAND_99;
  reg [63:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [63:0] _RAND_104;
  reg [63:0] _RAND_105;
  reg [63:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [63:0] _RAND_108;
  reg [63:0] _RAND_109;
  reg [63:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [63:0] _RAND_112;
  reg [63:0] _RAND_113;
  reg [63:0] _RAND_114;
  reg [63:0] _RAND_115;
  reg [63:0] _RAND_116;
  reg [63:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [63:0] _RAND_119;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [63:0] _RAND_123;
  reg [63:0] _RAND_124;
  reg [63:0] _RAND_125;
  reg [63:0] _RAND_126;
  reg [63:0] _RAND_127;
  reg [63:0] _RAND_128;
  reg [63:0] _RAND_129;
  reg [63:0] _RAND_130;
  reg [63:0] _RAND_131;
  reg [63:0] _RAND_132;
  reg [63:0] _RAND_133;
  reg [63:0] _RAND_134;
  reg [63:0] _RAND_135;
  reg [63:0] _RAND_136;
  reg [63:0] _RAND_137;
  reg [63:0] _RAND_138;
  reg [63:0] _RAND_139;
  reg [63:0] _RAND_140;
  reg [63:0] _RAND_141;
  reg [63:0] _RAND_142;
  reg [63:0] _RAND_143;
  reg [63:0] _RAND_144;
  reg [63:0] _RAND_145;
  reg [63:0] _RAND_146;
  reg [63:0] _RAND_147;
  reg [63:0] _RAND_148;
  reg [63:0] _RAND_149;
  reg [63:0] _RAND_150;
  reg [63:0] _RAND_151;
  reg [63:0] _RAND_152;
  reg [63:0] _RAND_153;
  reg [63:0] _RAND_154;
  reg [63:0] _RAND_155;
  reg [63:0] _RAND_156;
  reg [63:0] _RAND_157;
  reg [63:0] _RAND_158;
  reg [63:0] _RAND_159;
  reg [63:0] _RAND_160;
  reg [63:0] _RAND_161;
  reg [63:0] _RAND_162;
  reg [63:0] _RAND_163;
  reg [63:0] _RAND_164;
  reg [63:0] _RAND_165;
  reg [63:0] _RAND_166;
  reg [63:0] _RAND_167;
  reg [63:0] _RAND_168;
  reg [63:0] _RAND_169;
  reg [63:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [63:0] _RAND_172;
  reg [63:0] _RAND_173;
  reg [63:0] _RAND_174;
  reg [63:0] _RAND_175;
  reg [63:0] _RAND_176;
  reg [63:0] _RAND_177;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] mtvec; // @[CSR.scala 251:22]
  reg [63:0] mcounteren; // @[CSR.scala 252:27]
  reg [63:0] mcause; // @[CSR.scala 253:23]
  reg [63:0] mtval; // @[CSR.scala 254:22]
  reg [63:0] mepc; // @[CSR.scala 255:17]
  reg [63:0] mie; // @[CSR.scala 257:20]
  reg [63:0] mipReg; // @[CSR.scala 259:24]
  wire [11:0] _T_23 = {meip_0,1'h0,1'h0,1'h0,mtip_0,1'h0,2'h0,msip_0,3'h0}; // @[CSR.scala 261:22]
  wire [63:0] _GEN_331 = {{52'd0}, _T_23}; // @[CSR.scala 261:29]
  wire [63:0] _T_24 = _GEN_331 | mipReg; // @[CSR.scala 261:29]
  wire  mip_s_u = _T_24[0]; // @[CSR.scala 261:47]
  wire  mip_s_s = _T_24[1]; // @[CSR.scala 261:47]
  wire  mip_s_h = _T_24[2]; // @[CSR.scala 261:47]
  wire  mip_s_m = _T_24[3]; // @[CSR.scala 261:47]
  wire  mip_t_u = _T_24[4]; // @[CSR.scala 261:47]
  wire  mip_t_s = _T_24[5]; // @[CSR.scala 261:47]
  wire  mip_t_h = _T_24[6]; // @[CSR.scala 261:47]
  wire  mip_t_m = _T_24[7]; // @[CSR.scala 261:47]
  wire  mip_e_u = _T_24[8]; // @[CSR.scala 261:47]
  wire  mip_e_s = _T_24[9]; // @[CSR.scala 261:47]
  wire  mip_e_h = _T_24[10]; // @[CSR.scala 261:47]
  wire  mip_e_m = _T_24[11]; // @[CSR.scala 261:47]
  reg [63:0] misa; // @[CSR.scala 269:21]
  reg [63:0] mstatus; // @[CSR.scala 277:24]
  wire  mstatusStruct_ie_u = mstatus[0]; // @[CSR.scala 298:39]
  wire  mstatusStruct_ie_s = mstatus[1]; // @[CSR.scala 298:39]
  wire  mstatusStruct_ie_h = mstatus[2]; // @[CSR.scala 298:39]
  wire  mstatusStruct_ie_m = mstatus[3]; // @[CSR.scala 298:39]
  wire  mstatusStruct_pie_u = mstatus[4]; // @[CSR.scala 298:39]
  wire  mstatusStruct_pie_s = mstatus[5]; // @[CSR.scala 298:39]
  wire  mstatusStruct_pie_h = mstatus[6]; // @[CSR.scala 298:39]
  wire  mstatusStruct_pie_m = mstatus[7]; // @[CSR.scala 298:39]
  wire  mstatusStruct_spp = mstatus[8]; // @[CSR.scala 298:39]
  wire [1:0] mstatusStruct_hpp = mstatus[10:9]; // @[CSR.scala 298:39]
  wire [1:0] mstatusStruct_mpp = mstatus[12:11]; // @[CSR.scala 298:39]
  wire [1:0] mstatusStruct_fs = mstatus[14:13]; // @[CSR.scala 298:39]
  wire [1:0] mstatusStruct_xs = mstatus[16:15]; // @[CSR.scala 298:39]
  wire  mstatusStruct_mprv = mstatus[17]; // @[CSR.scala 298:39]
  wire  mstatusStruct_sum = mstatus[18]; // @[CSR.scala 298:39]
  wire  mstatusStruct_mxr = mstatus[19]; // @[CSR.scala 298:39]
  wire  mstatusStruct_tvm = mstatus[20]; // @[CSR.scala 298:39]
  wire  mstatusStruct_tw = mstatus[21]; // @[CSR.scala 298:39]
  wire  mstatusStruct_tsr = mstatus[22]; // @[CSR.scala 298:39]
  wire [8:0] mstatusStruct_pad0 = mstatus[31:23]; // @[CSR.scala 298:39]
  wire [1:0] mstatusStruct_uxl = mstatus[33:32]; // @[CSR.scala 298:39]
  wire [1:0] mstatusStruct_sxl = mstatus[35:34]; // @[CSR.scala 298:39]
  wire [26:0] mstatusStruct_pad1 = mstatus[62:36]; // @[CSR.scala 298:39]
  wire  mstatusStruct_sd = mstatus[63]; // @[CSR.scala 298:39]
  reg [63:0] medeleg; // @[CSR.scala 305:24]
  reg [63:0] mideleg; // @[CSR.scala 306:24]
  reg [63:0] mscratch; // @[CSR.scala 307:25]
  reg [63:0] pmpcfg0; // @[CSR.scala 309:24]
  reg [63:0] pmpcfg1; // @[CSR.scala 310:24]
  reg [63:0] pmpcfg2; // @[CSR.scala 311:24]
  reg [63:0] pmpcfg3; // @[CSR.scala 312:24]
  reg [63:0] pmpaddr0; // @[CSR.scala 313:25]
  reg [63:0] pmpaddr1; // @[CSR.scala 314:25]
  reg [63:0] pmpaddr2; // @[CSR.scala 315:25]
  reg [63:0] pmpaddr3; // @[CSR.scala 316:25]
  reg [63:0] stvec; // @[CSR.scala 330:22]
  wire [63:0] sieMask = 64'h222 & mideleg; // @[CSR.scala 332:26]
  reg [63:0] satp; // @[CSR.scala 335:21]
  reg [63:0] sepc; // @[CSR.scala 336:21]
  reg [63:0] scause; // @[CSR.scala 337:23]
  reg [63:0] stval; // @[CSR.scala 338:18]
  reg [63:0] sscratch; // @[CSR.scala 339:25]
  reg [63:0] scounteren; // @[CSR.scala 340:27]
  reg  lr; // @[CSR.scala 353:19]
  reg [63:0] lrAddr; // @[CSR.scala 354:23]
  reg [1:0] priviledgeMode; // @[CSR.scala 367:31]
  reg [63:0] perfCnts_0; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_1; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_2; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_3; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_4; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_5; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_6; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_7; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_8; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_9; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_10; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_11; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_12; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_13; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_14; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_15; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_16; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_17; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_18; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_19; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_20; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_21; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_22; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_23; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_24; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_25; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_26; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_27; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_28; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_29; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_30; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_31; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_32; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_33; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_34; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_35; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_36; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_37; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_38; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_39; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_40; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_41; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_42; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_43; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_44; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_45; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_46; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_47; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_48; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_49; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_50; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_51; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_52; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_53; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_54; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_55; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_56; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_57; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_58; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_59; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_60; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_61; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_62; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_63; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_64; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_65; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_66; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_67; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_68; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_69; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_70; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_71; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_72; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_73; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_74; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_75; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_76; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_77; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_78; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_79; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_80; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_81; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_82; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_83; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_84; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_85; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_86; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_87; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_88; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_89; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_90; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_91; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_92; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_93; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_94; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_95; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_96; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_97; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_98; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_99; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_100; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_101; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_102; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_103; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_104; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_105; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_106; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_107; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_108; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_109; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_110; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_111; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_112; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_113; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_114; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_115; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_116; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_117; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_118; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_119; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_120; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_121; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_122; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_123; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_124; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_125; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_126; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_127; // @[CSR.scala 372:47]
  wire [5:0] _T_732 = {mip_t_s,mip_t_u,mip_s_m,mip_s_h,mip_s_s,mip_s_u}; // @[CSR.scala 415:27]
  wire [11:0] _T_738 = {mip_e_m,mip_e_h,mip_e_s,mip_e_u,mip_t_m,mip_t_h,_T_732}; // @[CSR.scala 415:27]
  wire [11:0] addr = io_in_bits_src2[11:0]; // @[CSR.scala 455:18]
  wire [63:0] csri = {59'h0,io_cfIn_instr[19:15]}; // @[Cat.scala 29:58]
  wire  _T_1007 = 12'hb06 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1169 = _T_1007 ? perfCnts_6 : 64'h0; // @[Mux.scala 27:72]
  wire  _T_1008 = 12'hb49 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1170 = _T_1008 ? perfCnts_73 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1331 = _T_1169 | _T_1170; // @[Mux.scala 27:72]
  wire  _T_1009 = 12'hb3c == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1171 = _T_1009 ? perfCnts_60 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1332 = _T_1331 | _T_1171; // @[Mux.scala 27:72]
  wire  _T_1010 = 12'hb69 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1172 = _T_1010 ? perfCnts_105 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1333 = _T_1332 | _T_1172; // @[Mux.scala 27:72]
  wire  _T_1011 = 12'hb7c == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1173 = _T_1011 ? perfCnts_124 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1334 = _T_1333 | _T_1173; // @[Mux.scala 27:72]
  wire  _T_1012 = 12'hf12 == addr; // @[LookupTree.scala 24:34]
  wire  _T_1013 = 12'hb5c == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1175 = _T_1013 ? perfCnts_92 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1336 = _T_1334 | _T_1175; // @[Mux.scala 27:72]
  wire  _T_1014 = 12'hb15 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1176 = _T_1014 ? perfCnts_21 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1337 = _T_1336 | _T_1176; // @[Mux.scala 27:72]
  wire  _T_1015 = 12'hb26 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1177 = _T_1015 ? perfCnts_38 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1338 = _T_1337 | _T_1177; // @[Mux.scala 27:72]
  wire  _T_1016 = 12'h180 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1178 = _T_1016 ? satp : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1339 = _T_1338 | _T_1178; // @[Mux.scala 27:72]
  wire  _T_1017 = 12'hb66 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1179 = _T_1017 ? perfCnts_102 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1340 = _T_1339 | _T_1179; // @[Mux.scala 27:72]
  wire  _T_1018 = 12'hb75 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1180 = _T_1018 ? perfCnts_117 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1341 = _T_1340 | _T_1180; // @[Mux.scala 27:72]
  wire  _T_1019 = 12'hb55 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1181 = _T_1019 ? perfCnts_85 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1342 = _T_1341 | _T_1181; // @[Mux.scala 27:72]
  wire  _T_1020 = 12'h3b1 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1182 = _T_1020 ? pmpaddr1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1343 = _T_1342 | _T_1182; // @[Mux.scala 27:72]
  wire  _T_1021 = 12'hb1c == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1183 = _T_1021 ? perfCnts_28 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1344 = _T_1343 | _T_1183; // @[Mux.scala 27:72]
  wire  _T_1022 = 12'h3a2 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1184 = _T_1022 ? pmpcfg2 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1345 = _T_1344 | _T_1184; // @[Mux.scala 27:72]
  wire  _T_1023 = 12'hb46 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1185 = _T_1023 ? perfCnts_70 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1346 = _T_1345 | _T_1185; // @[Mux.scala 27:72]
  wire  _T_1024 = 12'h140 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1186 = _T_1024 ? sscratch : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1347 = _T_1346 | _T_1186; // @[Mux.scala 27:72]
  wire  _T_1025 = 12'hb09 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1187 = _T_1025 ? perfCnts_9 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1348 = _T_1347 | _T_1187; // @[Mux.scala 27:72]
  wire  _T_1026 = 12'hb03 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1188 = _T_1026 ? perfCnts_3 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1349 = _T_1348 | _T_1188; // @[Mux.scala 27:72]
  wire  _T_1027 = 12'hb35 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1189 = _T_1027 ? perfCnts_53 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1350 = _T_1349 | _T_1189; // @[Mux.scala 27:72]
  wire  _T_1028 = 12'hb64 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1190 = _T_1028 ? perfCnts_100 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1351 = _T_1350 | _T_1190; // @[Mux.scala 27:72]
  wire  _T_1029 = 12'hb51 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1191 = _T_1029 ? perfCnts_81 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1352 = _T_1351 | _T_1191; // @[Mux.scala 27:72]
  wire  _T_1030 = 12'hb29 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1192 = _T_1030 ? perfCnts_41 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1353 = _T_1352 | _T_1192; // @[Mux.scala 27:72]
  wire  _T_1031 = 12'h302 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1193 = _T_1031 ? medeleg : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1354 = _T_1353 | _T_1193; // @[Mux.scala 27:72]
  wire  _T_1032 = 12'hb71 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1194 = _T_1032 ? perfCnts_113 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1355 = _T_1354 | _T_1194; // @[Mux.scala 27:72]
  wire  _T_1033 = 12'hb24 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1195 = _T_1033 ? perfCnts_36 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1356 = _T_1355 | _T_1195; // @[Mux.scala 27:72]
  wire  _T_1034 = 12'h105 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1196 = _T_1034 ? stvec : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1357 = _T_1356 | _T_1196; // @[Mux.scala 27:72]
  wire  _T_1035 = 12'hb0d == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1197 = _T_1035 ? perfCnts_13 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1358 = _T_1357 | _T_1197; // @[Mux.scala 27:72]
  wire  _T_1036 = 12'hb4d == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1198 = _T_1036 ? perfCnts_77 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1359 = _T_1358 | _T_1198; // @[Mux.scala 27:72]
  wire  _T_1037 = 12'h141 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1199 = _T_1037 ? sepc : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1360 = _T_1359 | _T_1199; // @[Mux.scala 27:72]
  wire  _T_1038 = 12'hb40 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1200 = _T_1038 ? perfCnts_64 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1361 = _T_1360 | _T_1200; // @[Mux.scala 27:72]
  wire  _T_1039 = 12'h342 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1201 = _T_1039 ? mcause : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1362 = _T_1361 | _T_1201; // @[Mux.scala 27:72]
  wire  _T_1040 = 12'hb6d == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1202 = _T_1040 ? perfCnts_109 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1363 = _T_1362 | _T_1202; // @[Mux.scala 27:72]
  wire  _T_1041 = 12'hb11 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1203 = _T_1041 ? perfCnts_17 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1364 = _T_1363 | _T_1203; // @[Mux.scala 27:72]
  wire  _T_1042 = 12'hb2d == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1204 = _T_1042 ? perfCnts_45 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1365 = _T_1364 | _T_1204; // @[Mux.scala 27:72]
  wire  _T_1043 = 12'h306 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1205 = _T_1043 ? mcounteren : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1366 = _T_1365 | _T_1205; // @[Mux.scala 27:72]
  wire  _T_1044 = 12'hb44 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1206 = _T_1044 ? perfCnts_68 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1367 = _T_1366 | _T_1206; // @[Mux.scala 27:72]
  wire  _T_1045 = 12'hb6a == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1207 = _T_1045 ? perfCnts_106 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1368 = _T_1367 | _T_1207; // @[Mux.scala 27:72]
  wire  _T_1046 = 12'hf11 == addr; // @[LookupTree.scala 24:34]
  wire  _T_1047 = 12'hb5e == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1209 = _T_1047 ? perfCnts_94 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1370 = _T_1368 | _T_1209; // @[Mux.scala 27:72]
  wire  _T_1048 = 12'hb59 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1210 = _T_1048 ? perfCnts_89 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1371 = _T_1370 | _T_1210; // @[Mux.scala 27:72]
  wire  _T_1049 = 12'h104 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_887 = mie & sieMask; // @[RegMap.scala 48:84]
  wire [63:0] _T_1211 = _T_1049 ? _T_887 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1372 = _T_1371 | _T_1211; // @[Mux.scala 27:72]
  wire  _T_1050 = 12'hb79 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1212 = _T_1050 ? perfCnts_121 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1373 = _T_1372 | _T_1212; // @[Mux.scala 27:72]
  wire  _T_1051 = 12'hb4a == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1213 = _T_1051 ? perfCnts_74 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1374 = _T_1373 | _T_1213; // @[Mux.scala 27:72]
  wire  _T_1052 = 12'hb39 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1214 = _T_1052 ? perfCnts_57 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1375 = _T_1374 | _T_1214; // @[Mux.scala 27:72]
  wire  _T_1053 = 12'hb0a == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1215 = _T_1053 ? perfCnts_10 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1376 = _T_1375 | _T_1215; // @[Mux.scala 27:72]
  wire  _T_1054 = 12'hb04 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1216 = _T_1054 ? perfCnts_4 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1377 = _T_1376 | _T_1216; // @[Mux.scala 27:72]
  wire  _T_1055 = 12'hb38 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1217 = _T_1055 ? perfCnts_56 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1378 = _T_1377 | _T_1217; // @[Mux.scala 27:72]
  wire  _T_1056 = 12'h144 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _GEN_332 = {{52'd0}, _T_738}; // @[RegMap.scala 48:84]
  wire [63:0] _T_894 = _GEN_332 & sieMask; // @[RegMap.scala 48:84]
  wire [63:0] _T_1218 = _T_1056 ? _T_894 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1379 = _T_1378 | _T_1218; // @[Mux.scala 27:72]
  wire  _T_1057 = 12'hb18 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1219 = _T_1057 ? perfCnts_24 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1380 = _T_1379 | _T_1219; // @[Mux.scala 27:72]
  wire  _T_1058 = 12'hb4f == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1220 = _T_1058 ? perfCnts_79 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1381 = _T_1380 | _T_1220; // @[Mux.scala 27:72]
  wire  _T_1059 = 12'hb19 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1221 = _T_1059 ? perfCnts_25 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1382 = _T_1381 | _T_1221; // @[Mux.scala 27:72]
  wire  _T_1060 = 12'hb2a == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1222 = _T_1060 ? perfCnts_42 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1383 = _T_1382 | _T_1222; // @[Mux.scala 27:72]
  wire  _T_1061 = 12'h100 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_899 = mstatus & 64'h80000003000de122; // @[RegMap.scala 48:84]
  wire [63:0] _T_1223 = _T_1061 ? _T_899 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1384 = _T_1383 | _T_1223; // @[Mux.scala 27:72]
  wire  _T_1062 = 12'hb3d == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1224 = _T_1062 ? perfCnts_61 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1385 = _T_1384 | _T_1224; // @[Mux.scala 27:72]
  wire  _T_1063 = 12'hb0e == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1225 = _T_1063 ? perfCnts_14 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1386 = _T_1385 | _T_1225; // @[Mux.scala 27:72]
  wire  _T_1064 = 12'hb34 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1226 = _T_1064 ? perfCnts_52 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1387 = _T_1386 | _T_1226; // @[Mux.scala 27:72]
  wire  _T_1065 = 12'hb74 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1227 = _T_1065 ? perfCnts_116 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1388 = _T_1387 | _T_1227; // @[Mux.scala 27:72]
  wire  _T_1066 = 12'hb14 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1228 = _T_1066 ? perfCnts_20 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1389 = _T_1388 | _T_1228; // @[Mux.scala 27:72]
  wire  _T_1067 = 12'hb1d == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1229 = _T_1067 ? perfCnts_29 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1390 = _T_1389 | _T_1229; // @[Mux.scala 27:72]
  wire  _T_1068 = 12'hb54 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1230 = _T_1068 ? perfCnts_84 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1391 = _T_1390 | _T_1230; // @[Mux.scala 27:72]
  wire  _T_1069 = 12'hb23 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1231 = _T_1069 ? perfCnts_35 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1392 = _T_1391 | _T_1231; // @[Mux.scala 27:72]
  wire  _T_1070 = 12'hb2e == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1232 = _T_1070 ? perfCnts_46 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1393 = _T_1392 | _T_1232; // @[Mux.scala 27:72]
  wire  _T_1071 = 12'hb6e == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1233 = _T_1071 ? perfCnts_110 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1394 = _T_1393 | _T_1233; // @[Mux.scala 27:72]
  wire  _T_1072 = 12'hb43 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1234 = _T_1072 ? perfCnts_67 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1395 = _T_1394 | _T_1234; // @[Mux.scala 27:72]
  wire  _T_1073 = 12'hb63 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1235 = _T_1073 ? perfCnts_99 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1396 = _T_1395 | _T_1235; // @[Mux.scala 27:72]
  wire  _T_1074 = 12'h305 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1236 = _T_1074 ? mtvec : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1397 = _T_1396 | _T_1236; // @[Mux.scala 27:72]
  wire  _T_1075 = 12'hb5d == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1237 = _T_1075 ? perfCnts_93 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1398 = _T_1397 | _T_1237; // @[Mux.scala 27:72]
  wire  _T_1076 = 12'hb78 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1238 = _T_1076 ? perfCnts_120 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1399 = _T_1398 | _T_1238; // @[Mux.scala 27:72]
  wire  _T_1077 = 12'hb58 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1239 = _T_1077 ? perfCnts_88 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1400 = _T_1399 | _T_1239; // @[Mux.scala 27:72]
  wire  _T_1078 = 12'hb7d == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1240 = _T_1078 ? perfCnts_125 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1401 = _T_1400 | _T_1240; // @[Mux.scala 27:72]
  wire  _T_1079 = 12'hb4e == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1241 = _T_1079 ? perfCnts_78 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1402 = _T_1401 | _T_1241; // @[Mux.scala 27:72]
  wire  _T_1080 = 12'hb2b == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1242 = _T_1080 ? perfCnts_43 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1403 = _T_1402 | _T_1242; // @[Mux.scala 27:72]
  wire  _T_1081 = 12'hb7a == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1243 = _T_1081 ? perfCnts_122 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1404 = _T_1403 | _T_1243; // @[Mux.scala 27:72]
  wire  _T_1082 = 12'hb21 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1244 = _T_1082 ? perfCnts_33 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1405 = _T_1404 | _T_1244; // @[Mux.scala 27:72]
  wire  _T_1083 = 12'h304 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1245 = _T_1083 ? mie : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1406 = _T_1405 | _T_1245; // @[Mux.scala 27:72]
  wire  _T_1084 = 12'hb01 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1246 = _T_1084 ? perfCnts_1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1407 = _T_1406 | _T_1246; // @[Mux.scala 27:72]
  wire  _T_1085 = 12'hb0b == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1247 = _T_1085 ? perfCnts_11 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1408 = _T_1407 | _T_1247; // @[Mux.scala 27:72]
  wire  _T_1086 = 12'hb4b == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1248 = _T_1086 ? perfCnts_75 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1409 = _T_1408 | _T_1248; // @[Mux.scala 27:72]
  wire  _T_1087 = 12'hb77 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1249 = _T_1087 ? perfCnts_119 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1410 = _T_1409 | _T_1249; // @[Mux.scala 27:72]
  wire  _T_1088 = 12'h3b3 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1250 = _T_1088 ? pmpaddr3 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1411 = _T_1410 | _T_1250; // @[Mux.scala 27:72]
  wire  _T_1089 = 12'hb5a == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1251 = _T_1089 ? perfCnts_90 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1412 = _T_1411 | _T_1251; // @[Mux.scala 27:72]
  wire  _T_1090 = 12'hb17 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1252 = _T_1090 ? perfCnts_23 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1413 = _T_1412 | _T_1252; // @[Mux.scala 27:72]
  wire  _T_1091 = 12'hb7f == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1253 = _T_1091 ? perfCnts_127 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1414 = _T_1413 | _T_1253; // @[Mux.scala 27:72]
  wire  _T_1092 = 12'hb28 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1254 = _T_1092 ? perfCnts_40 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1415 = _T_1414 | _T_1254; // @[Mux.scala 27:72]
  wire  _T_1093 = 12'hb50 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1255 = _T_1093 ? perfCnts_80 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1416 = _T_1415 | _T_1255; // @[Mux.scala 27:72]
  wire  _T_1094 = 12'hb37 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1256 = _T_1094 ? perfCnts_55 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1417 = _T_1416 | _T_1256; // @[Mux.scala 27:72]
  wire  _T_1095 = 12'hb08 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1257 = _T_1095 ? perfCnts_8 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1418 = _T_1417 | _T_1257; // @[Mux.scala 27:72]
  wire  _T_1096 = 12'h143 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1258 = _T_1096 ? stval : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1419 = _T_1418 | _T_1258; // @[Mux.scala 27:72]
  wire  _T_1097 = 12'hb6b == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1259 = _T_1097 ? perfCnts_107 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1420 = _T_1419 | _T_1259; // @[Mux.scala 27:72]
  wire  _T_1098 = 12'hb3a == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1260 = _T_1098 ? perfCnts_58 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1421 = _T_1420 | _T_1260; // @[Mux.scala 27:72]
  wire  _T_1099 = 12'h301 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1261 = _T_1099 ? misa : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1422 = _T_1421 | _T_1261; // @[Mux.scala 27:72]
  wire  _T_1100 = 12'hb70 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1262 = _T_1100 ? perfCnts_112 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1423 = _T_1422 | _T_1262; // @[Mux.scala 27:72]
  wire  _T_1101 = 12'hb1a == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1263 = _T_1101 ? perfCnts_26 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1424 = _T_1423 | _T_1263; // @[Mux.scala 27:72]
  wire  _T_1102 = 12'hb5f == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1264 = _T_1102 ? perfCnts_95 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1425 = _T_1424 | _T_1264; // @[Mux.scala 27:72]
  wire  _T_1103 = 12'h300 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1265 = _T_1103 ? mstatus : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1426 = _T_1425 | _T_1265; // @[Mux.scala 27:72]
  wire  _T_1104 = 12'hb13 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1266 = _T_1104 ? perfCnts_19 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1427 = _T_1426 | _T_1266; // @[Mux.scala 27:72]
  wire  _T_1105 = 12'hb73 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1267 = _T_1105 ? perfCnts_115 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1428 = _T_1427 | _T_1267; // @[Mux.scala 27:72]
  wire  _T_1106 = 12'hb33 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1268 = _T_1106 ? perfCnts_51 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1429 = _T_1428 | _T_1268; // @[Mux.scala 27:72]
  wire  _T_1107 = 12'hb62 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1269 = _T_1107 ? perfCnts_98 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1430 = _T_1429 | _T_1269; // @[Mux.scala 27:72]
  wire  _T_1108 = 12'hb00 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1270 = _T_1108 ? perfCnts_0 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1431 = _T_1430 | _T_1270; // @[Mux.scala 27:72]
  wire  _T_1109 = 12'h3b0 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1271 = _T_1109 ? pmpaddr0 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1432 = _T_1431 | _T_1271; // @[Mux.scala 27:72]
  wire  _T_1110 = 12'hb3e == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1272 = _T_1110 ? perfCnts_62 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1433 = _T_1432 | _T_1272; // @[Mux.scala 27:72]
  wire  _T_1111 = 12'hb6f == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1273 = _T_1111 ? perfCnts_111 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1434 = _T_1433 | _T_1273; // @[Mux.scala 27:72]
  wire  _T_1112 = 12'hb1e == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1274 = _T_1112 ? perfCnts_30 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1435 = _T_1434 | _T_1274; // @[Mux.scala 27:72]
  wire  _T_1113 = 12'hb53 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1275 = _T_1113 ? perfCnts_83 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1436 = _T_1435 | _T_1275; // @[Mux.scala 27:72]
  wire  _T_1114 = 12'h344 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1276 = _T_1114 ? _GEN_332 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1437 = _T_1436 | _T_1276; // @[Mux.scala 27:72]
  wire  _T_1115 = 12'hb7e == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1277 = _T_1115 ? perfCnts_126 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1438 = _T_1437 | _T_1277; // @[Mux.scala 27:72]
  wire  _T_1116 = 12'hb2f == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1278 = _T_1116 ? perfCnts_47 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1439 = _T_1438 | _T_1278; // @[Mux.scala 27:72]
  wire  _T_1117 = 12'hb05 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1279 = _T_1117 ? perfCnts_5 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1440 = _T_1439 | _T_1279; // @[Mux.scala 27:72]
  wire  _T_1118 = 12'hb22 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1280 = _T_1118 ? perfCnts_34 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1441 = _T_1440 | _T_1280; // @[Mux.scala 27:72]
  wire  _T_1119 = 12'hb48 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1281 = _T_1119 ? perfCnts_72 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1442 = _T_1441 | _T_1281; // @[Mux.scala 27:72]
  wire  _T_1120 = 12'hb42 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1282 = _T_1120 ? perfCnts_66 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1443 = _T_1442 | _T_1282; // @[Mux.scala 27:72]
  wire  _T_1121 = 12'hb0f == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1283 = _T_1121 ? perfCnts_15 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1444 = _T_1443 | _T_1283; // @[Mux.scala 27:72]
  wire  _T_1122 = 12'hb68 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1284 = _T_1122 ? perfCnts_104 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1445 = _T_1444 | _T_1284; // @[Mux.scala 27:72]
  wire  _T_1123 = 12'hb57 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1285 = _T_1123 ? perfCnts_87 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1446 = _T_1445 | _T_1285; // @[Mux.scala 27:72]
  wire  _T_1124 = 12'hb16 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1286 = _T_1124 ? perfCnts_22 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1447 = _T_1446 | _T_1286; // @[Mux.scala 27:72]
  wire  _T_1125 = 12'hb1b == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1287 = _T_1125 ? perfCnts_27 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1448 = _T_1447 | _T_1287; // @[Mux.scala 27:72]
  wire  _T_1126 = 12'hb2c == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1288 = _T_1126 ? perfCnts_44 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1449 = _T_1448 | _T_1288; // @[Mux.scala 27:72]
  wire  _T_1127 = 12'hb7b == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1289 = _T_1127 ? perfCnts_123 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1450 = _T_1449 | _T_1289; // @[Mux.scala 27:72]
  wire  _T_1128 = 12'hb4c == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1290 = _T_1128 ? perfCnts_76 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1451 = _T_1450 | _T_1290; // @[Mux.scala 27:72]
  wire  _T_1129 = 12'hb20 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1291 = _T_1129 ? perfCnts_32 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1452 = _T_1451 | _T_1291; // @[Mux.scala 27:72]
  wire  _T_1130 = 12'hb31 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1292 = _T_1130 ? perfCnts_49 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1453 = _T_1452 | _T_1292; // @[Mux.scala 27:72]
  wire  _T_1131 = 12'hb3b == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1293 = _T_1131 ? perfCnts_59 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1454 = _T_1453 | _T_1293; // @[Mux.scala 27:72]
  wire  _T_1132 = 12'hb6c == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1294 = _T_1132 ? perfCnts_108 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1455 = _T_1454 | _T_1294; // @[Mux.scala 27:72]
  wire  _T_1133 = 12'hb02 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1295 = _T_1133 ? perfCnts_2 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1456 = _T_1455 | _T_1295; // @[Mux.scala 27:72]
  wire  _T_1134 = 12'h3a3 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1296 = _T_1134 ? pmpcfg3 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1457 = _T_1456 | _T_1296; // @[Mux.scala 27:72]
  wire  _T_1135 = 12'hb45 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1297 = _T_1135 ? perfCnts_69 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1458 = _T_1457 | _T_1297; // @[Mux.scala 27:72]
  wire  _T_1136 = 12'hb36 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1298 = _T_1136 ? perfCnts_54 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1459 = _T_1458 | _T_1298; // @[Mux.scala 27:72]
  wire  _T_1137 = 12'hb0c == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1299 = _T_1137 ? perfCnts_12 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1460 = _T_1459 | _T_1299; // @[Mux.scala 27:72]
  wire  _T_1138 = 12'hb67 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1300 = _T_1138 ? perfCnts_103 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1461 = _T_1460 | _T_1300; // @[Mux.scala 27:72]
  wire  _T_1139 = 12'h303 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1301 = _T_1139 ? mideleg : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1462 = _T_1461 | _T_1301; // @[Mux.scala 27:72]
  wire  _T_1140 = 12'hb5b == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1302 = _T_1140 ? perfCnts_91 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1463 = _T_1462 | _T_1302; // @[Mux.scala 27:72]
  wire  _T_1141 = 12'hb27 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1303 = _T_1141 ? perfCnts_39 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1464 = _T_1463 | _T_1303; // @[Mux.scala 27:72]
  wire  _T_1142 = 12'hb25 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1304 = _T_1142 ? perfCnts_37 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1465 = _T_1464 | _T_1304; // @[Mux.scala 27:72]
  wire  _T_1143 = 12'h3b2 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1305 = _T_1143 ? pmpaddr2 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1466 = _T_1465 | _T_1305; // @[Mux.scala 27:72]
  wire  _T_1144 = 12'hb07 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1306 = _T_1144 ? perfCnts_7 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1467 = _T_1466 | _T_1306; // @[Mux.scala 27:72]
  wire  _T_1145 = 12'hf13 == addr; // @[LookupTree.scala 24:34]
  wire  _T_1146 = 12'hb76 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1308 = _T_1146 ? perfCnts_118 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1469 = _T_1467 | _T_1308; // @[Mux.scala 27:72]
  wire  _T_1147 = 12'hb60 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1309 = _T_1147 ? perfCnts_96 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1470 = _T_1469 | _T_1309; // @[Mux.scala 27:72]
  wire  _T_1148 = 12'h3a1 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1310 = _T_1148 ? pmpcfg1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1471 = _T_1470 | _T_1310; // @[Mux.scala 27:72]
  wire  _T_1149 = 12'hb56 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1311 = _T_1149 ? perfCnts_86 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1472 = _T_1471 | _T_1311; // @[Mux.scala 27:72]
  wire  _T_1150 = 12'h340 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1312 = _T_1150 ? mscratch : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1473 = _T_1472 | _T_1312; // @[Mux.scala 27:72]
  wire  _T_1151 = 12'hb65 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1313 = _T_1151 ? perfCnts_101 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1474 = _T_1473 | _T_1313; // @[Mux.scala 27:72]
  wire  _T_1152 = 12'hb72 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1314 = _T_1152 ? perfCnts_114 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1475 = _T_1474 | _T_1314; // @[Mux.scala 27:72]
  wire  _T_1153 = 12'hf14 == addr; // @[LookupTree.scala 24:34]
  wire  _T_1154 = 12'h341 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1316 = _T_1154 ? mepc : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1477 = _T_1475 | _T_1316; // @[Mux.scala 27:72]
  wire  _T_1155 = 12'h343 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1317 = _T_1155 ? mtval : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1478 = _T_1477 | _T_1317; // @[Mux.scala 27:72]
  wire  _T_1156 = 12'h106 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1318 = _T_1156 ? scounteren : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1479 = _T_1478 | _T_1318; // @[Mux.scala 27:72]
  wire  _T_1157 = 12'hb61 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1319 = _T_1157 ? perfCnts_97 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1480 = _T_1479 | _T_1319; // @[Mux.scala 27:72]
  wire  _T_1158 = 12'h3a0 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1320 = _T_1158 ? pmpcfg0 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1481 = _T_1480 | _T_1320; // @[Mux.scala 27:72]
  wire  _T_1159 = 12'hb1f == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1321 = _T_1159 ? perfCnts_31 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1482 = _T_1481 | _T_1321; // @[Mux.scala 27:72]
  wire  _T_1160 = 12'hb52 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1322 = _T_1160 ? perfCnts_82 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1483 = _T_1482 | _T_1322; // @[Mux.scala 27:72]
  wire  _T_1161 = 12'hb30 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1323 = _T_1161 ? perfCnts_48 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1484 = _T_1483 | _T_1323; // @[Mux.scala 27:72]
  wire  _T_1162 = 12'h142 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1324 = _T_1162 ? scause : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1485 = _T_1484 | _T_1324; // @[Mux.scala 27:72]
  wire  _T_1163 = 12'hb3f == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1325 = _T_1163 ? perfCnts_63 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1486 = _T_1485 | _T_1325; // @[Mux.scala 27:72]
  wire  _T_1164 = 12'hb41 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1326 = _T_1164 ? perfCnts_65 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1487 = _T_1486 | _T_1326; // @[Mux.scala 27:72]
  wire  _T_1165 = 12'hb47 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1327 = _T_1165 ? perfCnts_71 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1488 = _T_1487 | _T_1327; // @[Mux.scala 27:72]
  wire  _T_1166 = 12'hb32 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1328 = _T_1166 ? perfCnts_50 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1489 = _T_1488 | _T_1328; // @[Mux.scala 27:72]
  wire  _T_1167 = 12'hb10 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1329 = _T_1167 ? perfCnts_16 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1490 = _T_1489 | _T_1329; // @[Mux.scala 27:72]
  wire  _T_1168 = 12'hb12 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1330 = _T_1168 ? perfCnts_18 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] rdata = _T_1490 | _T_1330; // @[Mux.scala 27:72]
  wire [63:0] _T_793 = rdata | io_in_bits_src1; // @[CSR.scala 460:30]
  wire [63:0] _T_794 = ~io_in_bits_src1; // @[CSR.scala 461:32]
  wire [63:0] _T_795 = rdata & _T_794; // @[CSR.scala 461:30]
  wire [63:0] _T_796 = rdata | csri; // @[CSR.scala 463:30]
  wire [63:0] _T_797 = ~csri; // @[CSR.scala 464:32]
  wire [63:0] _T_798 = rdata & _T_797; // @[CSR.scala 464:30]
  wire  _T_799 = 7'h1 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_800 = 7'h2 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_801 = 7'h3 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_802 = 7'h5 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_803 = 7'h6 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_804 = 7'h7 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire [63:0] _T_805 = _T_799 ? io_in_bits_src1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_806 = _T_800 ? _T_793 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_807 = _T_801 ? _T_795 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_808 = _T_802 ? csri : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_809 = _T_803 ? _T_796 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_810 = _T_804 ? _T_798 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_811 = _T_805 | _T_806; // @[Mux.scala 27:72]
  wire [63:0] _T_812 = _T_811 | _T_807; // @[Mux.scala 27:72]
  wire [63:0] _T_813 = _T_812 | _T_808; // @[Mux.scala 27:72]
  wire [63:0] _T_814 = _T_813 | _T_809; // @[Mux.scala 27:72]
  wire [63:0] wdata = _T_814 | _T_810; // @[Mux.scala 27:72]
  wire  _T_821 = wdata[63:60] == 4'h0; // @[CSR.scala 468:60]
  wire  _T_827 = wdata[63:60] == 4'h8; // @[CSR.scala 468:109]
  wire  satpLegalMode = _T_821 | _T_827; // @[CSR.scala 468:69]
  wire  _T_828 = io_in_bits_func != 7'h0; // @[CSR.scala 471:28]
  wire  _T_829 = io_in_valid & _T_828; // @[CSR.scala 471:20]
  wire  _T_830 = addr != 12'h180; // @[CSR.scala 471:56]
  wire  _T_831 = _T_830 | satpLegalMode; // @[CSR.scala 471:67]
  wire  wen = _T_829 & _T_831; // @[CSR.scala 471:47]
  wire  isIllegalMode = priviledgeMode < addr[9:8]; // @[CSR.scala 472:39]
  wire  _T_835 = io_in_bits_func == 7'h2; // @[CSR.scala 473:24]
  wire  _T_836 = io_in_bits_func == 7'h6; // @[CSR.scala 473:50]
  wire  _T_837 = _T_835 | _T_836; // @[CSR.scala 473:42]
  wire  _T_838 = io_in_bits_src1 == 64'h0; // @[CSR.scala 473:78]
  wire  justRead = _T_837 & _T_838; // @[CSR.scala 473:70]
  wire  _T_840 = addr[11:10] == 2'h3; // @[CSR.scala 474:45]
  wire  _T_841 = wen & _T_840; // @[CSR.scala 474:28]
  wire  _T_842 = ~justRead; // @[CSR.scala 474:61]
  wire  isIllegalWrite = _T_841 & _T_842; // @[CSR.scala 474:58]
  wire  isIllegalAccess = isIllegalMode | isIllegalWrite; // @[CSR.scala 475:39]
  wire  _T_843 = ~isIllegalAccess; // @[CSR.scala 477:54]
  wire  _T_844 = wen & _T_843; // @[CSR.scala 477:51]
  wire  _T_1493 = addr == 12'hb06; // @[RegMap.scala 50:65]
  wire  _T_1494 = _T_844 & _T_1493; // @[RegMap.scala 50:56]
  wire  _T_1499 = addr == 12'hb49; // @[RegMap.scala 50:65]
  wire  _T_1500 = _T_844 & _T_1499; // @[RegMap.scala 50:56]
  wire  _T_1505 = addr == 12'hb3c; // @[RegMap.scala 50:65]
  wire  _T_1506 = _T_844 & _T_1505; // @[RegMap.scala 50:56]
  wire  _T_1511 = addr == 12'hb69; // @[RegMap.scala 50:65]
  wire  _T_1512 = _T_844 & _T_1511; // @[RegMap.scala 50:56]
  wire  _T_1517 = addr == 12'hb7c; // @[RegMap.scala 50:65]
  wire  _T_1518 = _T_844 & _T_1517; // @[RegMap.scala 50:56]
  wire  _T_1523 = addr == 12'hb5c; // @[RegMap.scala 50:65]
  wire  _T_1524 = _T_844 & _T_1523; // @[RegMap.scala 50:56]
  wire  _T_1529 = addr == 12'hb15; // @[RegMap.scala 50:65]
  wire  _T_1530 = _T_844 & _T_1529; // @[RegMap.scala 50:56]
  wire  _T_1535 = addr == 12'hb26; // @[RegMap.scala 50:65]
  wire  _T_1536 = _T_844 & _T_1535; // @[RegMap.scala 50:56]
  wire  _T_1541 = addr == 12'h180; // @[RegMap.scala 50:65]
  wire  _T_1542 = _T_844 & _T_1541; // @[RegMap.scala 50:56]
  wire  _T_1547 = addr == 12'hb66; // @[RegMap.scala 50:65]
  wire  _T_1548 = _T_844 & _T_1547; // @[RegMap.scala 50:56]
  wire  _T_1553 = addr == 12'hb75; // @[RegMap.scala 50:65]
  wire  _T_1554 = _T_844 & _T_1553; // @[RegMap.scala 50:56]
  wire  _T_1559 = addr == 12'hb55; // @[RegMap.scala 50:65]
  wire  _T_1560 = _T_844 & _T_1559; // @[RegMap.scala 50:56]
  wire  _T_1565 = addr == 12'h3b1; // @[RegMap.scala 50:65]
  wire  _T_1566 = _T_844 & _T_1565; // @[RegMap.scala 50:56]
  wire  _T_1571 = addr == 12'hb1c; // @[RegMap.scala 50:65]
  wire  _T_1572 = _T_844 & _T_1571; // @[RegMap.scala 50:56]
  wire  _T_1577 = addr == 12'h3a2; // @[RegMap.scala 50:65]
  wire  _T_1578 = _T_844 & _T_1577; // @[RegMap.scala 50:56]
  wire  _T_1583 = addr == 12'hb46; // @[RegMap.scala 50:65]
  wire  _T_1584 = _T_844 & _T_1583; // @[RegMap.scala 50:56]
  wire  _T_1589 = addr == 12'h140; // @[RegMap.scala 50:65]
  wire  _T_1590 = _T_844 & _T_1589; // @[RegMap.scala 50:56]
  wire  _T_1595 = addr == 12'hb09; // @[RegMap.scala 50:65]
  wire  _T_1596 = _T_844 & _T_1595; // @[RegMap.scala 50:56]
  wire  _T_1601 = addr == 12'hb03; // @[RegMap.scala 50:65]
  wire  _T_1602 = _T_844 & _T_1601; // @[RegMap.scala 50:56]
  wire  _T_1607 = addr == 12'hb35; // @[RegMap.scala 50:65]
  wire  _T_1608 = _T_844 & _T_1607; // @[RegMap.scala 50:56]
  wire  _T_1619 = addr == 12'hb51; // @[RegMap.scala 50:65]
  wire  _T_1620 = _T_844 & _T_1619; // @[RegMap.scala 50:56]
  wire  _T_1625 = addr == 12'hb29; // @[RegMap.scala 50:65]
  wire  _T_1626 = _T_844 & _T_1625; // @[RegMap.scala 50:56]
  wire  _T_1631 = addr == 12'h302; // @[RegMap.scala 50:65]
  wire  _T_1632 = _T_844 & _T_1631; // @[RegMap.scala 50:56]
  wire [63:0] _T_1633 = wdata & 64'hbbff; // @[BitUtils.scala 32:13]
  wire [63:0] _T_1635 = medeleg & 64'h4400; // @[BitUtils.scala 32:36]
  wire [63:0] _T_1636 = _T_1633 | _T_1635; // @[BitUtils.scala 32:25]
  wire  _T_1637 = addr == 12'hb71; // @[RegMap.scala 50:65]
  wire  _T_1638 = _T_844 & _T_1637; // @[RegMap.scala 50:56]
  wire  _T_1643 = addr == 12'hb24; // @[RegMap.scala 50:65]
  wire  _T_1644 = _T_844 & _T_1643; // @[RegMap.scala 50:56]
  wire  _T_1649 = addr == 12'h105; // @[RegMap.scala 50:65]
  wire  _T_1650 = _T_844 & _T_1649; // @[RegMap.scala 50:56]
  wire  _T_1655 = addr == 12'hb0d; // @[RegMap.scala 50:65]
  wire  _T_1656 = _T_844 & _T_1655; // @[RegMap.scala 50:56]
  wire  _T_1661 = addr == 12'hb4d; // @[RegMap.scala 50:65]
  wire  _T_1662 = _T_844 & _T_1661; // @[RegMap.scala 50:56]
  wire  _T_1667 = addr == 12'h141; // @[RegMap.scala 50:65]
  wire  _T_1668 = _T_844 & _T_1667; // @[RegMap.scala 50:56]
  wire  _T_1673 = addr == 12'hb40; // @[RegMap.scala 50:65]
  wire  _T_1674 = _T_844 & _T_1673; // @[RegMap.scala 50:56]
  wire  _T_1679 = addr == 12'h342; // @[RegMap.scala 50:65]
  wire  _T_1680 = _T_844 & _T_1679; // @[RegMap.scala 50:56]
  wire  _T_1685 = addr == 12'hb6d; // @[RegMap.scala 50:65]
  wire  _T_1686 = _T_844 & _T_1685; // @[RegMap.scala 50:56]
  wire  _T_1691 = addr == 12'hb11; // @[RegMap.scala 50:65]
  wire  _T_1692 = _T_844 & _T_1691; // @[RegMap.scala 50:56]
  wire  _T_1697 = addr == 12'hb2d; // @[RegMap.scala 50:65]
  wire  _T_1698 = _T_844 & _T_1697; // @[RegMap.scala 50:56]
  wire  _T_1703 = addr == 12'h306; // @[RegMap.scala 50:65]
  wire  _T_1704 = _T_844 & _T_1703; // @[RegMap.scala 50:56]
  wire  _T_1709 = addr == 12'hb44; // @[RegMap.scala 50:65]
  wire  _T_1710 = _T_844 & _T_1709; // @[RegMap.scala 50:56]
  wire  _T_1715 = addr == 12'hb6a; // @[RegMap.scala 50:65]
  wire  _T_1716 = _T_844 & _T_1715; // @[RegMap.scala 50:56]
  wire  _T_1721 = addr == 12'hb5e; // @[RegMap.scala 50:65]
  wire  _T_1722 = _T_844 & _T_1721; // @[RegMap.scala 50:56]
  wire  _T_1727 = addr == 12'hb59; // @[RegMap.scala 50:65]
  wire  _T_1728 = _T_844 & _T_1727; // @[RegMap.scala 50:56]
  wire  _T_1733 = addr == 12'h104; // @[RegMap.scala 50:65]
  wire  _T_1734 = _T_844 & _T_1733; // @[RegMap.scala 50:56]
  wire [63:0] _T_1735 = wdata & sieMask; // @[BitUtils.scala 32:13]
  wire [63:0] _T_1736 = ~sieMask; // @[BitUtils.scala 32:38]
  wire [63:0] _T_1737 = mie & _T_1736; // @[BitUtils.scala 32:36]
  wire [63:0] _T_1738 = _T_1735 | _T_1737; // @[BitUtils.scala 32:25]
  wire  _T_1739 = addr == 12'hb79; // @[RegMap.scala 50:65]
  wire  _T_1740 = _T_844 & _T_1739; // @[RegMap.scala 50:56]
  wire  _T_1745 = addr == 12'hb4a; // @[RegMap.scala 50:65]
  wire  _T_1746 = _T_844 & _T_1745; // @[RegMap.scala 50:56]
  wire  _T_1751 = addr == 12'hb39; // @[RegMap.scala 50:65]
  wire  _T_1752 = _T_844 & _T_1751; // @[RegMap.scala 50:56]
  wire  _T_1757 = addr == 12'hb0a; // @[RegMap.scala 50:65]
  wire  _T_1758 = _T_844 & _T_1757; // @[RegMap.scala 50:56]
  wire  _T_1763 = addr == 12'hb04; // @[RegMap.scala 50:65]
  wire  _T_1764 = _T_844 & _T_1763; // @[RegMap.scala 50:56]
  wire  _T_1769 = addr == 12'hb38; // @[RegMap.scala 50:65]
  wire  _T_1770 = _T_844 & _T_1769; // @[RegMap.scala 50:56]
  wire  _T_1775 = addr == 12'hb18; // @[RegMap.scala 50:65]
  wire  _T_1776 = _T_844 & _T_1775; // @[RegMap.scala 50:56]
  wire  _T_1781 = addr == 12'hb4f; // @[RegMap.scala 50:65]
  wire  _T_1782 = _T_844 & _T_1781; // @[RegMap.scala 50:56]
  wire  _T_1787 = addr == 12'hb19; // @[RegMap.scala 50:65]
  wire  _T_1788 = _T_844 & _T_1787; // @[RegMap.scala 50:56]
  wire  _T_1793 = addr == 12'hb2a; // @[RegMap.scala 50:65]
  wire  _T_1794 = _T_844 & _T_1793; // @[RegMap.scala 50:56]
  wire  _T_1799 = addr == 12'h100; // @[RegMap.scala 50:65]
  wire  _T_1800 = _T_844 & _T_1799; // @[RegMap.scala 50:56]
  wire [63:0] _T_1801 = wdata & 64'hc6122; // @[BitUtils.scala 32:13]
  wire [63:0] _T_1803 = mstatus & 64'h39edd; // @[BitUtils.scala 32:36]
  wire [63:0] _T_1804 = _T_1801 | _T_1803; // @[BitUtils.scala 32:25]
  wire  _T_1832 = _T_1804[14:13] == 2'h3; // @[CSR.scala 301:40]
  wire [63:0] _T_1834 = {_T_1832,_T_1804[62:0]}; // @[Cat.scala 29:58]
  wire  _T_1835 = addr == 12'hb3d; // @[RegMap.scala 50:65]
  wire  _T_1836 = _T_844 & _T_1835; // @[RegMap.scala 50:56]
  wire  _T_1841 = addr == 12'hb0e; // @[RegMap.scala 50:65]
  wire  _T_1842 = _T_844 & _T_1841; // @[RegMap.scala 50:56]
  wire  _T_1847 = addr == 12'hb34; // @[RegMap.scala 50:65]
  wire  _T_1848 = _T_844 & _T_1847; // @[RegMap.scala 50:56]
  wire  _T_1853 = addr == 12'hb74; // @[RegMap.scala 50:65]
  wire  _T_1854 = _T_844 & _T_1853; // @[RegMap.scala 50:56]
  wire  _T_1859 = addr == 12'hb14; // @[RegMap.scala 50:65]
  wire  _T_1860 = _T_844 & _T_1859; // @[RegMap.scala 50:56]
  wire  _T_1865 = addr == 12'hb1d; // @[RegMap.scala 50:65]
  wire  _T_1866 = _T_844 & _T_1865; // @[RegMap.scala 50:56]
  wire  _T_1871 = addr == 12'hb54; // @[RegMap.scala 50:65]
  wire  _T_1872 = _T_844 & _T_1871; // @[RegMap.scala 50:56]
  wire  _T_1877 = addr == 12'hb23; // @[RegMap.scala 50:65]
  wire  _T_1878 = _T_844 & _T_1877; // @[RegMap.scala 50:56]
  wire  _T_1883 = addr == 12'hb2e; // @[RegMap.scala 50:65]
  wire  _T_1884 = _T_844 & _T_1883; // @[RegMap.scala 50:56]
  wire  _T_1889 = addr == 12'hb6e; // @[RegMap.scala 50:65]
  wire  _T_1890 = _T_844 & _T_1889; // @[RegMap.scala 50:56]
  wire  _T_1895 = addr == 12'hb43; // @[RegMap.scala 50:65]
  wire  _T_1896 = _T_844 & _T_1895; // @[RegMap.scala 50:56]
  wire  _T_1907 = addr == 12'h305; // @[RegMap.scala 50:65]
  wire  _T_1908 = _T_844 & _T_1907; // @[RegMap.scala 50:56]
  wire  _T_1913 = addr == 12'hb5d; // @[RegMap.scala 50:65]
  wire  _T_1914 = _T_844 & _T_1913; // @[RegMap.scala 50:56]
  wire  _T_1919 = addr == 12'hb78; // @[RegMap.scala 50:65]
  wire  _T_1920 = _T_844 & _T_1919; // @[RegMap.scala 50:56]
  wire  _T_1925 = addr == 12'hb58; // @[RegMap.scala 50:65]
  wire  _T_1926 = _T_844 & _T_1925; // @[RegMap.scala 50:56]
  wire  _T_1931 = addr == 12'hb7d; // @[RegMap.scala 50:65]
  wire  _T_1932 = _T_844 & _T_1931; // @[RegMap.scala 50:56]
  wire  _T_1937 = addr == 12'hb4e; // @[RegMap.scala 50:65]
  wire  _T_1938 = _T_844 & _T_1937; // @[RegMap.scala 50:56]
  wire  _T_1943 = addr == 12'hb2b; // @[RegMap.scala 50:65]
  wire  _T_1944 = _T_844 & _T_1943; // @[RegMap.scala 50:56]
  wire  _T_1949 = addr == 12'hb7a; // @[RegMap.scala 50:65]
  wire  _T_1950 = _T_844 & _T_1949; // @[RegMap.scala 50:56]
  wire  _T_1955 = addr == 12'hb21; // @[RegMap.scala 50:65]
  wire  _T_1956 = _T_844 & _T_1955; // @[RegMap.scala 50:56]
  wire  _T_1961 = addr == 12'h304; // @[RegMap.scala 50:65]
  wire  _T_1962 = _T_844 & _T_1961; // @[RegMap.scala 50:56]
  wire  _T_1967 = addr == 12'hb01; // @[RegMap.scala 50:65]
  wire  _T_1968 = _T_844 & _T_1967; // @[RegMap.scala 50:56]
  wire  _T_1973 = addr == 12'hb0b; // @[RegMap.scala 50:65]
  wire  _T_1974 = _T_844 & _T_1973; // @[RegMap.scala 50:56]
  wire  _T_1979 = addr == 12'hb4b; // @[RegMap.scala 50:65]
  wire  _T_1980 = _T_844 & _T_1979; // @[RegMap.scala 50:56]
  wire  _T_1985 = addr == 12'hb77; // @[RegMap.scala 50:65]
  wire  _T_1986 = _T_844 & _T_1985; // @[RegMap.scala 50:56]
  wire  _T_1991 = addr == 12'h3b3; // @[RegMap.scala 50:65]
  wire  _T_1992 = _T_844 & _T_1991; // @[RegMap.scala 50:56]
  wire  _T_1997 = addr == 12'hb5a; // @[RegMap.scala 50:65]
  wire  _T_1998 = _T_844 & _T_1997; // @[RegMap.scala 50:56]
  wire  _T_2003 = addr == 12'hb17; // @[RegMap.scala 50:65]
  wire  _T_2004 = _T_844 & _T_2003; // @[RegMap.scala 50:56]
  wire  _T_2009 = addr == 12'hb7f; // @[RegMap.scala 50:65]
  wire  _T_2010 = _T_844 & _T_2009; // @[RegMap.scala 50:56]
  wire  _T_2015 = addr == 12'hb28; // @[RegMap.scala 50:65]
  wire  _T_2016 = _T_844 & _T_2015; // @[RegMap.scala 50:56]
  wire  _T_2021 = addr == 12'hb50; // @[RegMap.scala 50:65]
  wire  _T_2022 = _T_844 & _T_2021; // @[RegMap.scala 50:56]
  wire  _T_2027 = addr == 12'hb37; // @[RegMap.scala 50:65]
  wire  _T_2028 = _T_844 & _T_2027; // @[RegMap.scala 50:56]
  wire  _T_2033 = addr == 12'hb08; // @[RegMap.scala 50:65]
  wire  _T_2034 = _T_844 & _T_2033; // @[RegMap.scala 50:56]
  wire  _T_2039 = addr == 12'h143; // @[RegMap.scala 50:65]
  wire  _T_2040 = _T_844 & _T_2039; // @[RegMap.scala 50:56]
  wire [63:0] _GEN_88 = _T_2040 ? wdata : stval; // @[RegMap.scala 50:72]
  wire  _T_2045 = addr == 12'hb6b; // @[RegMap.scala 50:65]
  wire  _T_2046 = _T_844 & _T_2045; // @[RegMap.scala 50:56]
  wire  _T_2051 = addr == 12'hb3a; // @[RegMap.scala 50:65]
  wire  _T_2052 = _T_844 & _T_2051; // @[RegMap.scala 50:56]
  wire  _T_2057 = addr == 12'h301; // @[RegMap.scala 50:65]
  wire  _T_2058 = _T_844 & _T_2057; // @[RegMap.scala 50:56]
  wire  _T_2063 = addr == 12'hb70; // @[RegMap.scala 50:65]
  wire  _T_2064 = _T_844 & _T_2063; // @[RegMap.scala 50:56]
  wire  _T_2069 = addr == 12'hb1a; // @[RegMap.scala 50:65]
  wire  _T_2070 = _T_844 & _T_2069; // @[RegMap.scala 50:56]
  wire  _T_2075 = addr == 12'hb5f; // @[RegMap.scala 50:65]
  wire  _T_2076 = _T_844 & _T_2075; // @[RegMap.scala 50:56]
  wire  _T_2081 = addr == 12'h300; // @[RegMap.scala 50:65]
  wire  _T_2082 = _T_844 & _T_2081; // @[RegMap.scala 50:56]
  wire  _T_2114 = wdata[14:13] == 2'h3; // @[CSR.scala 301:40]
  wire [63:0] _T_2116 = {_T_2114,wdata[62:0]}; // @[Cat.scala 29:58]
  wire  _T_2117 = addr == 12'hb13; // @[RegMap.scala 50:65]
  wire  _T_2118 = _T_844 & _T_2117; // @[RegMap.scala 50:56]
  wire  _T_2123 = addr == 12'hb73; // @[RegMap.scala 50:65]
  wire  _T_2124 = _T_844 & _T_2123; // @[RegMap.scala 50:56]
  wire  _T_2129 = addr == 12'hb33; // @[RegMap.scala 50:65]
  wire  _T_2130 = _T_844 & _T_2129; // @[RegMap.scala 50:56]
  wire  _T_2135 = addr == 12'hb62; // @[RegMap.scala 50:65]
  wire  _T_2136 = _T_844 & _T_2135; // @[RegMap.scala 50:56]
  wire  _T_2147 = addr == 12'h3b0; // @[RegMap.scala 50:65]
  wire  _T_2148 = _T_844 & _T_2147; // @[RegMap.scala 50:56]
  wire  _T_2153 = addr == 12'hb3e; // @[RegMap.scala 50:65]
  wire  _T_2154 = _T_844 & _T_2153; // @[RegMap.scala 50:56]
  wire  _T_2159 = addr == 12'hb6f; // @[RegMap.scala 50:65]
  wire  _T_2160 = _T_844 & _T_2159; // @[RegMap.scala 50:56]
  wire  _T_2165 = addr == 12'hb1e; // @[RegMap.scala 50:65]
  wire  _T_2166 = _T_844 & _T_2165; // @[RegMap.scala 50:56]
  wire  _T_2171 = addr == 12'hb53; // @[RegMap.scala 50:65]
  wire  _T_2172 = _T_844 & _T_2171; // @[RegMap.scala 50:56]
  wire  _T_2177 = addr == 12'hb7e; // @[RegMap.scala 50:65]
  wire  _T_2178 = _T_844 & _T_2177; // @[RegMap.scala 50:56]
  wire  _T_2183 = addr == 12'hb2f; // @[RegMap.scala 50:65]
  wire  _T_2184 = _T_844 & _T_2183; // @[RegMap.scala 50:56]
  wire  _T_2189 = addr == 12'hb05; // @[RegMap.scala 50:65]
  wire  _T_2190 = _T_844 & _T_2189; // @[RegMap.scala 50:56]
  wire  _T_2195 = addr == 12'hb22; // @[RegMap.scala 50:65]
  wire  _T_2196 = _T_844 & _T_2195; // @[RegMap.scala 50:56]
  wire  _T_2201 = addr == 12'hb48; // @[RegMap.scala 50:65]
  wire  _T_2202 = _T_844 & _T_2201; // @[RegMap.scala 50:56]
  wire  _T_2207 = addr == 12'hb42; // @[RegMap.scala 50:65]
  wire  _T_2208 = _T_844 & _T_2207; // @[RegMap.scala 50:56]
  wire  _T_2213 = addr == 12'hb0f; // @[RegMap.scala 50:65]
  wire  _T_2214 = _T_844 & _T_2213; // @[RegMap.scala 50:56]
  wire  _T_2219 = addr == 12'hb68; // @[RegMap.scala 50:65]
  wire  _T_2220 = _T_844 & _T_2219; // @[RegMap.scala 50:56]
  wire  _T_2225 = addr == 12'hb57; // @[RegMap.scala 50:65]
  wire  _T_2226 = _T_844 & _T_2225; // @[RegMap.scala 50:56]
  wire  _T_2231 = addr == 12'hb16; // @[RegMap.scala 50:65]
  wire  _T_2232 = _T_844 & _T_2231; // @[RegMap.scala 50:56]
  wire  _T_2237 = addr == 12'hb1b; // @[RegMap.scala 50:65]
  wire  _T_2238 = _T_844 & _T_2237; // @[RegMap.scala 50:56]
  wire  _T_2243 = addr == 12'hb2c; // @[RegMap.scala 50:65]
  wire  _T_2244 = _T_844 & _T_2243; // @[RegMap.scala 50:56]
  wire  _T_2249 = addr == 12'hb7b; // @[RegMap.scala 50:65]
  wire  _T_2250 = _T_844 & _T_2249; // @[RegMap.scala 50:56]
  wire  _T_2255 = addr == 12'hb4c; // @[RegMap.scala 50:65]
  wire  _T_2256 = _T_844 & _T_2255; // @[RegMap.scala 50:56]
  wire  _T_2261 = addr == 12'hb20; // @[RegMap.scala 50:65]
  wire  _T_2262 = _T_844 & _T_2261; // @[RegMap.scala 50:56]
  wire  _T_2267 = addr == 12'hb31; // @[RegMap.scala 50:65]
  wire  _T_2268 = _T_844 & _T_2267; // @[RegMap.scala 50:56]
  wire  _T_2273 = addr == 12'hb3b; // @[RegMap.scala 50:65]
  wire  _T_2274 = _T_844 & _T_2273; // @[RegMap.scala 50:56]
  wire  _T_2279 = addr == 12'hb6c; // @[RegMap.scala 50:65]
  wire  _T_2280 = _T_844 & _T_2279; // @[RegMap.scala 50:56]
  wire  _T_2285 = addr == 12'hb02; // @[RegMap.scala 50:65]
  wire  _T_2286 = _T_844 & _T_2285; // @[RegMap.scala 50:56]
  wire  _T_2291 = addr == 12'h3a3; // @[RegMap.scala 50:65]
  wire  _T_2292 = _T_844 & _T_2291; // @[RegMap.scala 50:56]
  wire  _T_2297 = addr == 12'hb45; // @[RegMap.scala 50:65]
  wire  _T_2298 = _T_844 & _T_2297; // @[RegMap.scala 50:56]
  wire  _T_2303 = addr == 12'hb36; // @[RegMap.scala 50:65]
  wire  _T_2304 = _T_844 & _T_2303; // @[RegMap.scala 50:56]
  wire  _T_2309 = addr == 12'hb0c; // @[RegMap.scala 50:65]
  wire  _T_2310 = _T_844 & _T_2309; // @[RegMap.scala 50:56]
  wire  _T_2315 = addr == 12'hb67; // @[RegMap.scala 50:65]
  wire  _T_2316 = _T_844 & _T_2315; // @[RegMap.scala 50:56]
  wire  _T_2321 = addr == 12'h303; // @[RegMap.scala 50:65]
  wire  _T_2322 = _T_844 & _T_2321; // @[RegMap.scala 50:56]
  wire [63:0] _T_2323 = wdata & 64'h222; // @[BitUtils.scala 32:13]
  wire [63:0] _T_2325 = mideleg & 64'h1dd; // @[BitUtils.scala 32:36]
  wire [63:0] _T_2326 = _T_2323 | _T_2325; // @[BitUtils.scala 32:25]
  wire  _T_2327 = addr == 12'hb5b; // @[RegMap.scala 50:65]
  wire  _T_2328 = _T_844 & _T_2327; // @[RegMap.scala 50:56]
  wire  _T_2333 = addr == 12'hb27; // @[RegMap.scala 50:65]
  wire  _T_2334 = _T_844 & _T_2333; // @[RegMap.scala 50:56]
  wire  _T_2339 = addr == 12'hb25; // @[RegMap.scala 50:65]
  wire  _T_2340 = _T_844 & _T_2339; // @[RegMap.scala 50:56]
  wire  _T_2345 = addr == 12'h3b2; // @[RegMap.scala 50:65]
  wire  _T_2346 = _T_844 & _T_2345; // @[RegMap.scala 50:56]
  wire  _T_2351 = addr == 12'hb07; // @[RegMap.scala 50:65]
  wire  _T_2352 = _T_844 & _T_2351; // @[RegMap.scala 50:56]
  wire  _T_2357 = addr == 12'hb76; // @[RegMap.scala 50:65]
  wire  _T_2358 = _T_844 & _T_2357; // @[RegMap.scala 50:56]
  wire  _T_2363 = addr == 12'hb60; // @[RegMap.scala 50:65]
  wire  _T_2364 = _T_844 & _T_2363; // @[RegMap.scala 50:56]
  wire  _T_2369 = addr == 12'h3a1; // @[RegMap.scala 50:65]
  wire  _T_2370 = _T_844 & _T_2369; // @[RegMap.scala 50:56]
  wire  _T_2375 = addr == 12'hb56; // @[RegMap.scala 50:65]
  wire  _T_2376 = _T_844 & _T_2375; // @[RegMap.scala 50:56]
  wire  _T_2381 = addr == 12'h340; // @[RegMap.scala 50:65]
  wire  _T_2382 = _T_844 & _T_2381; // @[RegMap.scala 50:56]
  wire  _T_2393 = addr == 12'hb72; // @[RegMap.scala 50:65]
  wire  _T_2394 = _T_844 & _T_2393; // @[RegMap.scala 50:56]
  wire  _T_2399 = addr == 12'h341; // @[RegMap.scala 50:65]
  wire  _T_2400 = _T_844 & _T_2399; // @[RegMap.scala 50:56]
  wire  _T_2405 = addr == 12'h343; // @[RegMap.scala 50:65]
  wire  _T_2406 = _T_844 & _T_2405; // @[RegMap.scala 50:56]
  wire [63:0] _GEN_144 = _T_2406 ? wdata : mtval; // @[RegMap.scala 50:72]
  wire  _T_2411 = addr == 12'h106; // @[RegMap.scala 50:65]
  wire  _T_2412 = _T_844 & _T_2411; // @[RegMap.scala 50:56]
  wire  _T_2417 = addr == 12'hb61; // @[RegMap.scala 50:65]
  wire  _T_2418 = _T_844 & _T_2417; // @[RegMap.scala 50:56]
  wire  _T_2423 = addr == 12'h3a0; // @[RegMap.scala 50:65]
  wire  _T_2424 = _T_844 & _T_2423; // @[RegMap.scala 50:56]
  wire  _T_2429 = addr == 12'hb1f; // @[RegMap.scala 50:65]
  wire  _T_2430 = _T_844 & _T_2429; // @[RegMap.scala 50:56]
  wire  _T_2435 = addr == 12'hb52; // @[RegMap.scala 50:65]
  wire  _T_2436 = _T_844 & _T_2435; // @[RegMap.scala 50:56]
  wire  _T_2441 = addr == 12'hb30; // @[RegMap.scala 50:65]
  wire  _T_2442 = _T_844 & _T_2441; // @[RegMap.scala 50:56]
  wire  _T_2447 = addr == 12'h142; // @[RegMap.scala 50:65]
  wire  _T_2448 = _T_844 & _T_2447; // @[RegMap.scala 50:56]
  wire  _T_2453 = addr == 12'hb3f; // @[RegMap.scala 50:65]
  wire  _T_2454 = _T_844 & _T_2453; // @[RegMap.scala 50:56]
  wire  _T_2459 = addr == 12'hb41; // @[RegMap.scala 50:65]
  wire  _T_2460 = _T_844 & _T_2459; // @[RegMap.scala 50:56]
  wire  _T_2465 = addr == 12'hb47; // @[RegMap.scala 50:65]
  wire  _T_2466 = _T_844 & _T_2465; // @[RegMap.scala 50:56]
  wire  _T_2471 = addr == 12'hb32; // @[RegMap.scala 50:65]
  wire  _T_2472 = _T_844 & _T_2471; // @[RegMap.scala 50:56]
  wire  _T_2477 = addr == 12'hb10; // @[RegMap.scala 50:65]
  wire  _T_2478 = _T_844 & _T_2477; // @[RegMap.scala 50:56]
  wire  _T_2483 = addr == 12'hb12; // @[RegMap.scala 50:65]
  wire  _T_2484 = _T_844 & _T_2483; // @[RegMap.scala 50:56]
  wire  _T_2490 = _T_1007 ? 1'h0 : 1'h1; // @[Mux.scala 80:57]
  wire  _T_2492 = _T_1008 ? 1'h0 : _T_2490; // @[Mux.scala 80:57]
  wire  _T_2494 = _T_1009 ? 1'h0 : _T_2492; // @[Mux.scala 80:57]
  wire  _T_2496 = _T_1010 ? 1'h0 : _T_2494; // @[Mux.scala 80:57]
  wire  _T_2498 = _T_1011 ? 1'h0 : _T_2496; // @[Mux.scala 80:57]
  wire  _T_2500 = _T_1012 ? 1'h0 : _T_2498; // @[Mux.scala 80:57]
  wire  _T_2502 = _T_1013 ? 1'h0 : _T_2500; // @[Mux.scala 80:57]
  wire  _T_2504 = _T_1014 ? 1'h0 : _T_2502; // @[Mux.scala 80:57]
  wire  _T_2506 = _T_1015 ? 1'h0 : _T_2504; // @[Mux.scala 80:57]
  wire  _T_2508 = _T_1016 ? 1'h0 : _T_2506; // @[Mux.scala 80:57]
  wire  _T_2510 = _T_1017 ? 1'h0 : _T_2508; // @[Mux.scala 80:57]
  wire  _T_2512 = _T_1018 ? 1'h0 : _T_2510; // @[Mux.scala 80:57]
  wire  _T_2514 = _T_1019 ? 1'h0 : _T_2512; // @[Mux.scala 80:57]
  wire  _T_2516 = _T_1020 ? 1'h0 : _T_2514; // @[Mux.scala 80:57]
  wire  _T_2518 = _T_1021 ? 1'h0 : _T_2516; // @[Mux.scala 80:57]
  wire  _T_2520 = _T_1022 ? 1'h0 : _T_2518; // @[Mux.scala 80:57]
  wire  _T_2522 = _T_1023 ? 1'h0 : _T_2520; // @[Mux.scala 80:57]
  wire  _T_2524 = _T_1024 ? 1'h0 : _T_2522; // @[Mux.scala 80:57]
  wire  _T_2526 = _T_1025 ? 1'h0 : _T_2524; // @[Mux.scala 80:57]
  wire  _T_2528 = _T_1026 ? 1'h0 : _T_2526; // @[Mux.scala 80:57]
  wire  _T_2530 = _T_1027 ? 1'h0 : _T_2528; // @[Mux.scala 80:57]
  wire  _T_2532 = _T_1028 ? 1'h0 : _T_2530; // @[Mux.scala 80:57]
  wire  _T_2534 = _T_1029 ? 1'h0 : _T_2532; // @[Mux.scala 80:57]
  wire  _T_2536 = _T_1030 ? 1'h0 : _T_2534; // @[Mux.scala 80:57]
  wire  _T_2538 = _T_1031 ? 1'h0 : _T_2536; // @[Mux.scala 80:57]
  wire  _T_2540 = _T_1032 ? 1'h0 : _T_2538; // @[Mux.scala 80:57]
  wire  _T_2542 = _T_1033 ? 1'h0 : _T_2540; // @[Mux.scala 80:57]
  wire  _T_2544 = _T_1034 ? 1'h0 : _T_2542; // @[Mux.scala 80:57]
  wire  _T_2546 = _T_1035 ? 1'h0 : _T_2544; // @[Mux.scala 80:57]
  wire  _T_2548 = _T_1036 ? 1'h0 : _T_2546; // @[Mux.scala 80:57]
  wire  _T_2550 = _T_1037 ? 1'h0 : _T_2548; // @[Mux.scala 80:57]
  wire  _T_2552 = _T_1038 ? 1'h0 : _T_2550; // @[Mux.scala 80:57]
  wire  _T_2554 = _T_1039 ? 1'h0 : _T_2552; // @[Mux.scala 80:57]
  wire  _T_2556 = _T_1040 ? 1'h0 : _T_2554; // @[Mux.scala 80:57]
  wire  _T_2558 = _T_1041 ? 1'h0 : _T_2556; // @[Mux.scala 80:57]
  wire  _T_2560 = _T_1042 ? 1'h0 : _T_2558; // @[Mux.scala 80:57]
  wire  _T_2562 = _T_1043 ? 1'h0 : _T_2560; // @[Mux.scala 80:57]
  wire  _T_2564 = _T_1044 ? 1'h0 : _T_2562; // @[Mux.scala 80:57]
  wire  _T_2566 = _T_1045 ? 1'h0 : _T_2564; // @[Mux.scala 80:57]
  wire  _T_2568 = _T_1046 ? 1'h0 : _T_2566; // @[Mux.scala 80:57]
  wire  _T_2570 = _T_1047 ? 1'h0 : _T_2568; // @[Mux.scala 80:57]
  wire  _T_2572 = _T_1048 ? 1'h0 : _T_2570; // @[Mux.scala 80:57]
  wire  _T_2574 = _T_1049 ? 1'h0 : _T_2572; // @[Mux.scala 80:57]
  wire  _T_2576 = _T_1050 ? 1'h0 : _T_2574; // @[Mux.scala 80:57]
  wire  _T_2578 = _T_1051 ? 1'h0 : _T_2576; // @[Mux.scala 80:57]
  wire  _T_2580 = _T_1052 ? 1'h0 : _T_2578; // @[Mux.scala 80:57]
  wire  _T_2582 = _T_1053 ? 1'h0 : _T_2580; // @[Mux.scala 80:57]
  wire  _T_2584 = _T_1054 ? 1'h0 : _T_2582; // @[Mux.scala 80:57]
  wire  _T_2586 = _T_1055 ? 1'h0 : _T_2584; // @[Mux.scala 80:57]
  wire  _T_2588 = _T_1056 ? 1'h0 : _T_2586; // @[Mux.scala 80:57]
  wire  _T_2590 = _T_1057 ? 1'h0 : _T_2588; // @[Mux.scala 80:57]
  wire  _T_2592 = _T_1058 ? 1'h0 : _T_2590; // @[Mux.scala 80:57]
  wire  _T_2594 = _T_1059 ? 1'h0 : _T_2592; // @[Mux.scala 80:57]
  wire  _T_2596 = _T_1060 ? 1'h0 : _T_2594; // @[Mux.scala 80:57]
  wire  _T_2598 = _T_1061 ? 1'h0 : _T_2596; // @[Mux.scala 80:57]
  wire  _T_2600 = _T_1062 ? 1'h0 : _T_2598; // @[Mux.scala 80:57]
  wire  _T_2602 = _T_1063 ? 1'h0 : _T_2600; // @[Mux.scala 80:57]
  wire  _T_2604 = _T_1064 ? 1'h0 : _T_2602; // @[Mux.scala 80:57]
  wire  _T_2606 = _T_1065 ? 1'h0 : _T_2604; // @[Mux.scala 80:57]
  wire  _T_2608 = _T_1066 ? 1'h0 : _T_2606; // @[Mux.scala 80:57]
  wire  _T_2610 = _T_1067 ? 1'h0 : _T_2608; // @[Mux.scala 80:57]
  wire  _T_2612 = _T_1068 ? 1'h0 : _T_2610; // @[Mux.scala 80:57]
  wire  _T_2614 = _T_1069 ? 1'h0 : _T_2612; // @[Mux.scala 80:57]
  wire  _T_2616 = _T_1070 ? 1'h0 : _T_2614; // @[Mux.scala 80:57]
  wire  _T_2618 = _T_1071 ? 1'h0 : _T_2616; // @[Mux.scala 80:57]
  wire  _T_2620 = _T_1072 ? 1'h0 : _T_2618; // @[Mux.scala 80:57]
  wire  _T_2622 = _T_1073 ? 1'h0 : _T_2620; // @[Mux.scala 80:57]
  wire  _T_2624 = _T_1074 ? 1'h0 : _T_2622; // @[Mux.scala 80:57]
  wire  _T_2626 = _T_1075 ? 1'h0 : _T_2624; // @[Mux.scala 80:57]
  wire  _T_2628 = _T_1076 ? 1'h0 : _T_2626; // @[Mux.scala 80:57]
  wire  _T_2630 = _T_1077 ? 1'h0 : _T_2628; // @[Mux.scala 80:57]
  wire  _T_2632 = _T_1078 ? 1'h0 : _T_2630; // @[Mux.scala 80:57]
  wire  _T_2634 = _T_1079 ? 1'h0 : _T_2632; // @[Mux.scala 80:57]
  wire  _T_2636 = _T_1080 ? 1'h0 : _T_2634; // @[Mux.scala 80:57]
  wire  _T_2638 = _T_1081 ? 1'h0 : _T_2636; // @[Mux.scala 80:57]
  wire  _T_2640 = _T_1082 ? 1'h0 : _T_2638; // @[Mux.scala 80:57]
  wire  _T_2642 = _T_1083 ? 1'h0 : _T_2640; // @[Mux.scala 80:57]
  wire  _T_2644 = _T_1084 ? 1'h0 : _T_2642; // @[Mux.scala 80:57]
  wire  _T_2646 = _T_1085 ? 1'h0 : _T_2644; // @[Mux.scala 80:57]
  wire  _T_2648 = _T_1086 ? 1'h0 : _T_2646; // @[Mux.scala 80:57]
  wire  _T_2650 = _T_1087 ? 1'h0 : _T_2648; // @[Mux.scala 80:57]
  wire  _T_2652 = _T_1088 ? 1'h0 : _T_2650; // @[Mux.scala 80:57]
  wire  _T_2654 = _T_1089 ? 1'h0 : _T_2652; // @[Mux.scala 80:57]
  wire  _T_2656 = _T_1090 ? 1'h0 : _T_2654; // @[Mux.scala 80:57]
  wire  _T_2658 = _T_1091 ? 1'h0 : _T_2656; // @[Mux.scala 80:57]
  wire  _T_2660 = _T_1092 ? 1'h0 : _T_2658; // @[Mux.scala 80:57]
  wire  _T_2662 = _T_1093 ? 1'h0 : _T_2660; // @[Mux.scala 80:57]
  wire  _T_2664 = _T_1094 ? 1'h0 : _T_2662; // @[Mux.scala 80:57]
  wire  _T_2666 = _T_1095 ? 1'h0 : _T_2664; // @[Mux.scala 80:57]
  wire  _T_2668 = _T_1096 ? 1'h0 : _T_2666; // @[Mux.scala 80:57]
  wire  _T_2670 = _T_1097 ? 1'h0 : _T_2668; // @[Mux.scala 80:57]
  wire  _T_2672 = _T_1098 ? 1'h0 : _T_2670; // @[Mux.scala 80:57]
  wire  _T_2674 = _T_1099 ? 1'h0 : _T_2672; // @[Mux.scala 80:57]
  wire  _T_2676 = _T_1100 ? 1'h0 : _T_2674; // @[Mux.scala 80:57]
  wire  _T_2678 = _T_1101 ? 1'h0 : _T_2676; // @[Mux.scala 80:57]
  wire  _T_2680 = _T_1102 ? 1'h0 : _T_2678; // @[Mux.scala 80:57]
  wire  _T_2682 = _T_1103 ? 1'h0 : _T_2680; // @[Mux.scala 80:57]
  wire  _T_2684 = _T_1104 ? 1'h0 : _T_2682; // @[Mux.scala 80:57]
  wire  _T_2686 = _T_1105 ? 1'h0 : _T_2684; // @[Mux.scala 80:57]
  wire  _T_2688 = _T_1106 ? 1'h0 : _T_2686; // @[Mux.scala 80:57]
  wire  _T_2690 = _T_1107 ? 1'h0 : _T_2688; // @[Mux.scala 80:57]
  wire  _T_2692 = _T_1108 ? 1'h0 : _T_2690; // @[Mux.scala 80:57]
  wire  _T_2694 = _T_1109 ? 1'h0 : _T_2692; // @[Mux.scala 80:57]
  wire  _T_2696 = _T_1110 ? 1'h0 : _T_2694; // @[Mux.scala 80:57]
  wire  _T_2698 = _T_1111 ? 1'h0 : _T_2696; // @[Mux.scala 80:57]
  wire  _T_2700 = _T_1112 ? 1'h0 : _T_2698; // @[Mux.scala 80:57]
  wire  _T_2702 = _T_1113 ? 1'h0 : _T_2700; // @[Mux.scala 80:57]
  wire  _T_2704 = _T_1114 ? 1'h0 : _T_2702; // @[Mux.scala 80:57]
  wire  _T_2706 = _T_1115 ? 1'h0 : _T_2704; // @[Mux.scala 80:57]
  wire  _T_2708 = _T_1116 ? 1'h0 : _T_2706; // @[Mux.scala 80:57]
  wire  _T_2710 = _T_1117 ? 1'h0 : _T_2708; // @[Mux.scala 80:57]
  wire  _T_2712 = _T_1118 ? 1'h0 : _T_2710; // @[Mux.scala 80:57]
  wire  _T_2714 = _T_1119 ? 1'h0 : _T_2712; // @[Mux.scala 80:57]
  wire  _T_2716 = _T_1120 ? 1'h0 : _T_2714; // @[Mux.scala 80:57]
  wire  _T_2718 = _T_1121 ? 1'h0 : _T_2716; // @[Mux.scala 80:57]
  wire  _T_2720 = _T_1122 ? 1'h0 : _T_2718; // @[Mux.scala 80:57]
  wire  _T_2722 = _T_1123 ? 1'h0 : _T_2720; // @[Mux.scala 80:57]
  wire  _T_2724 = _T_1124 ? 1'h0 : _T_2722; // @[Mux.scala 80:57]
  wire  _T_2726 = _T_1125 ? 1'h0 : _T_2724; // @[Mux.scala 80:57]
  wire  _T_2728 = _T_1126 ? 1'h0 : _T_2726; // @[Mux.scala 80:57]
  wire  _T_2730 = _T_1127 ? 1'h0 : _T_2728; // @[Mux.scala 80:57]
  wire  _T_2732 = _T_1128 ? 1'h0 : _T_2730; // @[Mux.scala 80:57]
  wire  _T_2734 = _T_1129 ? 1'h0 : _T_2732; // @[Mux.scala 80:57]
  wire  _T_2736 = _T_1130 ? 1'h0 : _T_2734; // @[Mux.scala 80:57]
  wire  _T_2738 = _T_1131 ? 1'h0 : _T_2736; // @[Mux.scala 80:57]
  wire  _T_2740 = _T_1132 ? 1'h0 : _T_2738; // @[Mux.scala 80:57]
  wire  _T_2742 = _T_1133 ? 1'h0 : _T_2740; // @[Mux.scala 80:57]
  wire  _T_2744 = _T_1134 ? 1'h0 : _T_2742; // @[Mux.scala 80:57]
  wire  _T_2746 = _T_1135 ? 1'h0 : _T_2744; // @[Mux.scala 80:57]
  wire  _T_2748 = _T_1136 ? 1'h0 : _T_2746; // @[Mux.scala 80:57]
  wire  _T_2750 = _T_1137 ? 1'h0 : _T_2748; // @[Mux.scala 80:57]
  wire  _T_2752 = _T_1138 ? 1'h0 : _T_2750; // @[Mux.scala 80:57]
  wire  _T_2754 = _T_1139 ? 1'h0 : _T_2752; // @[Mux.scala 80:57]
  wire  _T_2756 = _T_1140 ? 1'h0 : _T_2754; // @[Mux.scala 80:57]
  wire  _T_2758 = _T_1141 ? 1'h0 : _T_2756; // @[Mux.scala 80:57]
  wire  _T_2760 = _T_1142 ? 1'h0 : _T_2758; // @[Mux.scala 80:57]
  wire  _T_2762 = _T_1143 ? 1'h0 : _T_2760; // @[Mux.scala 80:57]
  wire  _T_2764 = _T_1144 ? 1'h0 : _T_2762; // @[Mux.scala 80:57]
  wire  _T_2766 = _T_1145 ? 1'h0 : _T_2764; // @[Mux.scala 80:57]
  wire  _T_2768 = _T_1146 ? 1'h0 : _T_2766; // @[Mux.scala 80:57]
  wire  _T_2770 = _T_1147 ? 1'h0 : _T_2768; // @[Mux.scala 80:57]
  wire  _T_2772 = _T_1148 ? 1'h0 : _T_2770; // @[Mux.scala 80:57]
  wire  _T_2774 = _T_1149 ? 1'h0 : _T_2772; // @[Mux.scala 80:57]
  wire  _T_2776 = _T_1150 ? 1'h0 : _T_2774; // @[Mux.scala 80:57]
  wire  _T_2778 = _T_1151 ? 1'h0 : _T_2776; // @[Mux.scala 80:57]
  wire  _T_2780 = _T_1152 ? 1'h0 : _T_2778; // @[Mux.scala 80:57]
  wire  _T_2782 = _T_1153 ? 1'h0 : _T_2780; // @[Mux.scala 80:57]
  wire  _T_2784 = _T_1154 ? 1'h0 : _T_2782; // @[Mux.scala 80:57]
  wire  _T_2786 = _T_1155 ? 1'h0 : _T_2784; // @[Mux.scala 80:57]
  wire  _T_2788 = _T_1156 ? 1'h0 : _T_2786; // @[Mux.scala 80:57]
  wire  _T_2790 = _T_1157 ? 1'h0 : _T_2788; // @[Mux.scala 80:57]
  wire  _T_2792 = _T_1158 ? 1'h0 : _T_2790; // @[Mux.scala 80:57]
  wire  _T_2794 = _T_1159 ? 1'h0 : _T_2792; // @[Mux.scala 80:57]
  wire  _T_2796 = _T_1160 ? 1'h0 : _T_2794; // @[Mux.scala 80:57]
  wire  _T_2798 = _T_1161 ? 1'h0 : _T_2796; // @[Mux.scala 80:57]
  wire  _T_2800 = _T_1162 ? 1'h0 : _T_2798; // @[Mux.scala 80:57]
  wire  _T_2802 = _T_1163 ? 1'h0 : _T_2800; // @[Mux.scala 80:57]
  wire  _T_2804 = _T_1164 ? 1'h0 : _T_2802; // @[Mux.scala 80:57]
  wire  _T_2806 = _T_1165 ? 1'h0 : _T_2804; // @[Mux.scala 80:57]
  wire  _T_2808 = _T_1166 ? 1'h0 : _T_2806; // @[Mux.scala 80:57]
  wire  _T_2810 = _T_1167 ? 1'h0 : _T_2808; // @[Mux.scala 80:57]
  wire  isIllegalAddr = _T_1168 ? 1'h0 : _T_2810; // @[Mux.scala 80:57]
  wire  resetSatp = _T_1541 & wen; // @[CSR.scala 479:35]
  wire  _T_2825 = addr == 12'h344; // @[RegMap.scala 50:65]
  wire  _T_2826 = _T_844 & _T_2825; // @[RegMap.scala 50:56]
  wire [63:0] _T_2827 = wdata & 64'h77f; // @[BitUtils.scala 32:13]
  wire [63:0] _T_2829 = mipReg & 64'h80; // @[BitUtils.scala 32:36]
  wire [63:0] _T_2830 = _T_2827 | _T_2829; // @[BitUtils.scala 32:25]
  wire  _T_2831 = addr == 12'h144; // @[RegMap.scala 50:65]
  wire  _T_2832 = _T_844 & _T_2831; // @[RegMap.scala 50:56]
  wire [63:0] _T_2835 = mipReg & _T_1736; // @[BitUtils.scala 32:36]
  wire [63:0] _T_2836 = _T_1735 | _T_2835; // @[BitUtils.scala 32:25]
  wire  _T_2837 = addr == 12'h1; // @[CSR.scala 492:23]
  wire  _T_2838 = io_in_bits_func == 7'h0; // @[CSR.scala 492:46]
  wire  isEbreak = _T_2837 & _T_2838; // @[CSR.scala 492:38]
  wire  _T_2841 = addr == 12'h0; // @[CSR.scala 493:22]
  wire  isEcall = _T_2841 & _T_2838; // @[CSR.scala 493:36]
  wire  isMret = _T_1631 & _T_2838; // @[CSR.scala 494:36]
  wire  _T_2849 = addr == 12'h102; // @[CSR.scala 495:21]
  wire  isSret = _T_2849 & _T_2838; // @[CSR.scala 495:36]
  wire  _T_2853 = addr == 12'h2; // @[CSR.scala 496:21]
  wire  isUret = _T_2853 & _T_2838; // @[CSR.scala 496:36]
  reg [63:0] _T_2857; // @[GTimer.scala 24:20]
  wire [63:0] _T_2859 = _T_2857 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_2861 = wen & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  wire  _T_2863 = ~reset; // @[Debug.scala 56:24]
  reg [63:0] _T_2866; // @[GTimer.scala 24:20]
  wire [63:0] _T_2868 = _T_2866 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_2869; // @[GTimer.scala 24:20]
  wire [63:0] _T_2871 = _T_2869 + 64'h1; // @[GTimer.scala 25:12]
  wire  hasInstrPageFault = io_cfIn_exceptionVec_12 & io_in_valid; // @[CSR.scala 553:63]
  wire  _T_2884 = hasInstrPageFault | io_dmemMMU_loadPF; // @[CSR.scala 562:26]
  wire  _T_2885 = _T_2884 | io_dmemMMU_storePF; // @[CSR.scala 562:46]
  wire [38:0] _T_2887 = io_cfIn_pc + 39'h2; // @[CSR.scala 563:88]
  wire [24:0] _T_2891 = _T_2887[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_2892 = {_T_2891,_T_2887}; // @[Cat.scala 29:58]
  wire [24:0] _T_2896 = io_cfIn_pc[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_2897 = {_T_2896,io_cfIn_pc}; // @[Cat.scala 29:58]
  wire [63:0] _T_2898 = io_cfIn_crossPageIPFFix ? _T_2892 : _T_2897; // @[CSR.scala 563:42]
  wire [24:0] _T_2901 = io_dmemMMU_addr[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_2902 = {_T_2901,io_dmemMMU_addr}; // @[Cat.scala 29:58]
  wire [63:0] _T_2903 = hasInstrPageFault ? _T_2898 : _T_2902; // @[CSR.scala 563:19]
  wire  _T_2904 = priviledgeMode == 2'h3; // @[CSR.scala 564:25]
  reg [63:0] _T_2905; // @[GTimer.scala 24:20]
  wire [63:0] _T_2907 = _T_2905 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_2912; // @[GTimer.scala 24:20]
  wire [63:0] _T_2914 = _T_2912 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_2921 = io_cfIn_exceptionVec_4 | io_cfIn_exceptionVec_6; // @[CSR.scala 572:30]
  wire [38:0] dmemAddrMisalignedAddr = LSUADDR[38:0]; // @[CSR.scala 541:36 CSR.scala 559:28]
  wire [24:0] _T_2924 = dmemAddrMisalignedAddr[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_2925 = {_T_2924,dmemAddrMisalignedAddr}; // @[Cat.scala 29:58]
  reg [63:0] _T_2926; // @[GTimer.scala 24:20]
  wire [63:0] _T_2928 = _T_2926 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_2933; // @[GTimer.scala 24:20]
  wire [63:0] _T_2935 = _T_2933 + 64'h1; // @[GTimer.scala 25:12]
  wire  mipRaiseIntr_e_s = mip_e_s | meip_0; // @[CSR.scala 596:31]
  wire [11:0] _T_2953 = {mip_e_m,mip_e_h,mipRaiseIntr_e_s,mip_e_u,mip_t_m,mip_t_h,_T_732}; // @[CSR.scala 598:41]
  wire [63:0] _GEN_333 = {{52'd0}, _T_2953}; // @[CSR.scala 598:26]
  wire [63:0] ideleg = mideleg & _GEN_333; // @[CSR.scala 598:26]
  wire  _T_3018 = priviledgeMode == 2'h1; // @[CSR.scala 599:72]
  wire  _T_3019 = _T_3018 & mstatusStruct_ie_s; // @[CSR.scala 599:83]
  wire  _T_3020 = priviledgeMode < 2'h1; // @[CSR.scala 599:125]
  wire  _T_3021 = _T_3019 | _T_3020; // @[CSR.scala 599:106]
  wire  _T_3023 = _T_2904 & mstatusStruct_ie_m; // @[CSR.scala 600:64]
  wire  _T_3024 = priviledgeMode < 2'h3; // @[CSR.scala 600:106]
  wire  _T_3025 = _T_3023 | _T_3024; // @[CSR.scala 600:87]
  wire  intrVecEnable_0 = ideleg[0] ? _T_3021 : _T_3025; // @[CSR.scala 599:51]
  wire  intrVecEnable_1 = ideleg[1] ? _T_3021 : _T_3025; // @[CSR.scala 599:51]
  wire  intrVecEnable_2 = ideleg[2] ? _T_3021 : _T_3025; // @[CSR.scala 599:51]
  wire  intrVecEnable_3 = ideleg[3] ? _T_3021 : _T_3025; // @[CSR.scala 599:51]
  wire  intrVecEnable_4 = ideleg[4] ? _T_3021 : _T_3025; // @[CSR.scala 599:51]
  wire  intrVecEnable_5 = ideleg[5] ? _T_3021 : _T_3025; // @[CSR.scala 599:51]
  wire  intrVecEnable_6 = ideleg[6] ? _T_3021 : _T_3025; // @[CSR.scala 599:51]
  wire  intrVecEnable_7 = ideleg[7] ? _T_3021 : _T_3025; // @[CSR.scala 599:51]
  wire  intrVecEnable_8 = ideleg[8] ? _T_3021 : _T_3025; // @[CSR.scala 599:51]
  wire  intrVecEnable_9 = ideleg[9] ? _T_3021 : _T_3025; // @[CSR.scala 599:51]
  wire  intrVecEnable_10 = ideleg[10] ? _T_3021 : _T_3025; // @[CSR.scala 599:51]
  wire  intrVecEnable_11 = ideleg[11] ? _T_3021 : _T_3025; // @[CSR.scala 599:51]
  wire [11:0] _T_3138 = mie[11:0] & _T_2953; // @[CSR.scala 604:27]
  wire [5:0] _T_3143 = {intrVecEnable_5,intrVecEnable_4,intrVecEnable_3,intrVecEnable_2,intrVecEnable_1,intrVecEnable_0}; // @[CSR.scala 604:65]
  wire [11:0] _T_3149 = {intrVecEnable_11,intrVecEnable_10,intrVecEnable_9,intrVecEnable_8,intrVecEnable_7,intrVecEnable_6,_T_3143}; // @[CSR.scala 604:65]
  wire [11:0] intrVec = _T_3138 & _T_3149; // @[CSR.scala 604:49]
  wire [2:0] _T_3150 = io_cfIn_intrVec_4 ? 3'h4 : 3'h0; // @[CSR.scala 608:69]
  wire [3:0] _T_3151 = io_cfIn_intrVec_8 ? 4'h8 : {{1'd0}, _T_3150}; // @[CSR.scala 608:69]
  wire [3:0] _T_3152 = io_cfIn_intrVec_0 ? 4'h0 : _T_3151; // @[CSR.scala 608:69]
  wire [3:0] _T_3153 = io_cfIn_intrVec_5 ? 4'h5 : _T_3152; // @[CSR.scala 608:69]
  wire [3:0] _T_3154 = io_cfIn_intrVec_9 ? 4'h9 : _T_3153; // @[CSR.scala 608:69]
  wire [3:0] _T_3155 = io_cfIn_intrVec_1 ? 4'h1 : _T_3154; // @[CSR.scala 608:69]
  wire [3:0] _T_3156 = io_cfIn_intrVec_7 ? 4'h7 : _T_3155; // @[CSR.scala 608:69]
  wire [3:0] _T_3157 = io_cfIn_intrVec_11 ? 4'hb : _T_3156; // @[CSR.scala 608:69]
  wire [3:0] intrNO = io_cfIn_intrVec_3 ? 4'h3 : _T_3157; // @[CSR.scala 608:69]
  wire [5:0] _T_3162 = {io_cfIn_intrVec_5,io_cfIn_intrVec_4,io_cfIn_intrVec_3,io_cfIn_intrVec_2,io_cfIn_intrVec_1,io_cfIn_intrVec_0}; // @[CSR.scala 610:35]
  wire [11:0] _T_3168 = {io_cfIn_intrVec_11,io_cfIn_intrVec_10,io_cfIn_intrVec_9,io_cfIn_intrVec_8,io_cfIn_intrVec_7,io_cfIn_intrVec_6,_T_3162}; // @[CSR.scala 610:35]
  wire  raiseIntr = |_T_3168; // @[CSR.scala 610:42]
  wire  csrExceptionVec_3 = io_in_valid & isEbreak; // @[CSR.scala 617:46]
  wire  _T_3171 = _T_2904 & io_in_valid; // @[CSR.scala 618:55]
  wire  csrExceptionVec_11 = _T_3171 & isEcall; // @[CSR.scala 618:70]
  wire  _T_3174 = _T_3018 & io_in_valid; // @[CSR.scala 619:55]
  wire  csrExceptionVec_9 = _T_3174 & isEcall; // @[CSR.scala 619:70]
  wire  _T_3176 = priviledgeMode == 2'h0; // @[CSR.scala 620:45]
  wire  _T_3177 = _T_3176 & io_in_valid; // @[CSR.scala 620:55]
  wire  csrExceptionVec_8 = _T_3177 & isEcall; // @[CSR.scala 620:70]
  wire  _T_3179 = isIllegalAddr | isIllegalAccess; // @[CSR.scala 621:51]
  wire  csrExceptionVec_2 = _T_3179 & wen; // @[CSR.scala 621:71]
  wire [7:0] _T_3189 = {4'h0,csrExceptionVec_3,csrExceptionVec_2,2'h0}; // @[CSR.scala 625:49]
  wire [15:0] _T_3197 = {io_dmemMMU_storePF,1'h0,io_dmemMMU_loadPF,1'h0,csrExceptionVec_11,1'h0,csrExceptionVec_9,csrExceptionVec_8,_T_3189}; // @[CSR.scala 625:49]
  wire [7:0] _T_3204 = {1'h0,io_cfIn_exceptionVec_6,1'h0,io_cfIn_exceptionVec_4,1'h0,io_cfIn_exceptionVec_2,io_cfIn_exceptionVec_1,1'h0}; // @[CSR.scala 625:76]
  wire [15:0] _T_3212 = {2'h0,1'h0,io_cfIn_exceptionVec_12,4'h0,_T_3204}; // @[CSR.scala 625:76]
  wire [15:0] raiseExceptionVec = _T_3197 | _T_3212; // @[CSR.scala 625:52]
  wire  raiseException = |raiseExceptionVec; // @[CSR.scala 626:42]
  wire [2:0] _T_3214 = raiseExceptionVec[5] ? 3'h5 : 3'h0; // @[CSR.scala 627:74]
  wire [2:0] _T_3216 = raiseExceptionVec[7] ? 3'h7 : _T_3214; // @[CSR.scala 627:74]
  wire [3:0] _T_3218 = raiseExceptionVec[13] ? 4'hd : {{1'd0}, _T_3216}; // @[CSR.scala 627:74]
  wire [3:0] _T_3220 = raiseExceptionVec[15] ? 4'hf : _T_3218; // @[CSR.scala 627:74]
  wire [3:0] _T_3222 = raiseExceptionVec[4] ? 4'h4 : _T_3220; // @[CSR.scala 627:74]
  wire [3:0] _T_3224 = raiseExceptionVec[6] ? 4'h6 : _T_3222; // @[CSR.scala 627:74]
  wire [3:0] _T_3226 = raiseExceptionVec[8] ? 4'h8 : _T_3224; // @[CSR.scala 627:74]
  wire [3:0] _T_3228 = raiseExceptionVec[9] ? 4'h9 : _T_3226; // @[CSR.scala 627:74]
  wire [3:0] _T_3230 = raiseExceptionVec[11] ? 4'hb : _T_3228; // @[CSR.scala 627:74]
  wire [3:0] _T_3232 = raiseExceptionVec[0] ? 4'h0 : _T_3230; // @[CSR.scala 627:74]
  wire [3:0] _T_3234 = raiseExceptionVec[2] ? 4'h2 : _T_3232; // @[CSR.scala 627:74]
  wire [3:0] _T_3236 = raiseExceptionVec[1] ? 4'h1 : _T_3234; // @[CSR.scala 627:74]
  wire [3:0] _T_3238 = raiseExceptionVec[12] ? 4'hc : _T_3236; // @[CSR.scala 627:74]
  wire [3:0] exceptionNO = raiseExceptionVec[3] ? 4'h3 : _T_3238; // @[CSR.scala 627:74]
  wire [63:0] _T_3240 = {raiseIntr, 63'h0}; // @[CSR.scala 630:28]
  wire [3:0] _T_3241 = raiseIntr ? intrNO : exceptionNO; // @[CSR.scala 630:46]
  wire [63:0] _GEN_334 = {{60'd0}, _T_3241}; // @[CSR.scala 630:41]
  wire [63:0] causeNO = _T_3240 | _GEN_334; // @[CSR.scala 630:41]
  wire  _T_3243 = raiseException | raiseIntr; // @[CSR.scala 633:44]
  wire  raiseExceptionIntr = _T_3243 & io_instrValid; // @[CSR.scala 633:58]
  wire  _T_3245 = io_in_valid & _T_2838; // @[CSR.scala 636:31]
  wire  _T_3246 = _T_3245 | raiseExceptionIntr; // @[CSR.scala 636:58]
  wire [38:0] _T_3249 = io_cfIn_pc + 39'h4; // @[CSR.scala 638:51]
  wire [63:0] deleg = raiseIntr ? mideleg : medeleg; // @[CSR.scala 648:18]
  wire [63:0] _T_3342 = deleg >> causeNO[3:0]; // @[CSR.scala 650:22]
  wire  delegS = _T_3342[0] & _T_3024; // @[CSR.scala 650:38]
  wire [63:0] _T_3352 = delegS ? stvec : mtvec; // @[CSR.scala 654:20]
  wire [38:0] trapTarget = _T_3352[38:0]; // @[CSR.scala 654:42]
  wire  _T_3513 = io_in_valid & isUret; // @[CSR.scala 685:15]
  wire  _T_3433 = io_in_valid & isSret; // @[CSR.scala 672:15]
  wire  _T_3354 = io_in_valid & isMret; // @[CSR.scala 659:15]
  wire [38:0] _GEN_172 = _T_3433 ? sepc[38:0] : mepc[38:0]; // @[CSR.scala 672:26]
  wire [38:0] retTarget = _T_3513 ? 39'h0 : _GEN_172; // @[CSR.scala 685:26]
  wire [38:0] _T_3250 = raiseExceptionIntr ? trapTarget : retTarget; // @[CSR.scala 638:61]
  reg [63:0] _T_3282; // @[GTimer.scala 24:20]
  wire [63:0] _T_3284 = _T_3282 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_3286 = raiseExceptionIntr & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  reg [63:0] _T_3302; // @[GTimer.scala 24:20]
  wire [63:0] _T_3304 = _T_3302 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_3311; // @[GTimer.scala 24:20]
  wire [63:0] _T_3313 = _T_3311 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_3314; // @[GTimer.scala 24:20]
  wire [63:0] _T_3316 = _T_3314 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_3323; // @[GTimer.scala 24:20]
  wire [63:0] _T_3325 = _T_3323 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_3327 = io_redirect_valid & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  reg [63:0] _T_3332; // @[GTimer.scala 24:20]
  wire [63:0] _T_3334 = _T_3332 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_3336 = resetSatp & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  wire  _T_3347 = _T_2885 | io_cfIn_exceptionVec_4; // @[CSR.scala 651:78]
  wire  _T_3348 = _T_3347 | io_cfIn_exceptionVec_6; // @[CSR.scala 651:103]
  wire  _T_3349 = ~_T_3348; // @[CSR.scala 651:17]
  wire  tvalWen = _T_3349 | raiseIntr; // @[CSR.scala 651:130]
  wire [5:0] _T_3413 = {mstatusStruct_pie_s,mstatusStruct_pie_u,mstatusStruct_pie_m,mstatusStruct_ie_h,mstatusStruct_ie_s,mstatusStruct_ie_u}; // @[CSR.scala 667:27]
  wire [14:0] _T_3419 = {mstatusStruct_fs,2'h0,mstatusStruct_hpp,mstatusStruct_spp,1'h1,mstatusStruct_pie_h,_T_3413}; // @[CSR.scala 667:27]
  wire [6:0] _T_3424 = {mstatusStruct_tw,mstatusStruct_tvm,mstatusStruct_mxr,mstatusStruct_sum,mstatusStruct_mprv,mstatusStruct_xs}; // @[CSR.scala 667:27]
  wire [63:0] _T_3431 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,mstatusStruct_pad0,mstatusStruct_tsr,_T_3424,_T_3419}; // @[CSR.scala 667:27]
  wire [1:0] _T_3488 = {1'h0,mstatusStruct_spp}; // @[Cat.scala 29:58]
  wire [5:0] _T_3493 = {1'h1,mstatusStruct_pie_u,mstatusStruct_ie_m,mstatusStruct_ie_h,mstatusStruct_pie_s,mstatusStruct_ie_u}; // @[CSR.scala 680:27]
  wire [14:0] _T_3499 = {mstatusStruct_fs,mstatusStruct_mpp,mstatusStruct_hpp,1'h0,mstatusStruct_pie_m,mstatusStruct_pie_h,_T_3493}; // @[CSR.scala 680:27]
  wire [63:0] _T_3511 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,mstatusStruct_pad0,mstatusStruct_tsr,_T_3424,_T_3499}; // @[CSR.scala 680:27]
  wire [5:0] _T_3572 = {mstatusStruct_pie_s,1'h1,mstatusStruct_ie_m,mstatusStruct_ie_h,mstatusStruct_ie_s,mstatusStruct_pie_u}; // @[CSR.scala 692:27]
  wire [14:0] _T_3578 = {mstatusStruct_fs,mstatusStruct_mpp,mstatusStruct_hpp,mstatusStruct_spp,mstatusStruct_pie_m,mstatusStruct_pie_h,_T_3572}; // @[CSR.scala 692:27]
  wire [63:0] _T_3590 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,mstatusStruct_pad0,mstatusStruct_tsr,_T_3424,_T_3578}; // @[CSR.scala 692:27]
  wire [1:0] _GEN_180 = delegS ? priviledgeMode : {{1'd0}, mstatusStruct_spp}; // @[CSR.scala 700:19]
  wire  _GEN_181 = delegS ? mstatusStruct_ie_s : mstatusStruct_pie_s; // @[CSR.scala 700:19]
  wire  _GEN_182 = delegS ? 1'h0 : mstatusStruct_ie_s; // @[CSR.scala 700:19]
  wire [1:0] _GEN_187 = delegS ? mstatusStruct_mpp : priviledgeMode; // @[CSR.scala 700:19]
  wire  _GEN_188 = delegS ? mstatusStruct_pie_m : mstatusStruct_ie_m; // @[CSR.scala 700:19]
  wire  _GEN_189 = delegS & mstatusStruct_ie_m; // @[CSR.scala 700:19]
  wire [5:0] _T_3658 = {_GEN_181,mstatusStruct_pie_u,_GEN_189,mstatusStruct_ie_h,_GEN_182,mstatusStruct_ie_u}; // @[CSR.scala 727:27]
  wire [14:0] _T_3664 = {mstatusStruct_fs,_GEN_187,mstatusStruct_hpp,_GEN_180[0],_GEN_188,mstatusStruct_pie_h,_T_3658}; // @[CSR.scala 727:27]
  wire [63:0] _T_3676 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,mstatusStruct_pad0,mstatusStruct_tsr,_T_3424,_T_3664}; // @[CSR.scala 727:27]
  wire [63:0] _T_3678 = perfCnts_0 + 64'h1; // @[CSR.scala 837:71]
  wire  _T_3941 = 1'h1;
  wire [63:0] _T_3682 = perfCnts_2 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3684 = perfCnts_3 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3686 = perfCnts_4 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3688 = perfCnts_5 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3690 = perfCnts_6 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3692 = perfCnts_7 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3694 = perfCnts_8 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3696 = perfCnts_9 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3698 = perfCnts_10 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3700 = perfCnts_11 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3706 = perfCnts_14 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3708 = perfCnts_15 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3710 = perfCnts_16 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3712 = perfCnts_17 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3714 = perfCnts_18 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3716 = perfCnts_19 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3718 = perfCnts_20 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3720 = perfCnts_21 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3722 = perfCnts_22 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3724 = perfCnts_23 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3728 = perfCnts_25 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3730 = perfCnts_26 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3732 = perfCnts_27 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3734 = perfCnts_28 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3736 = perfCnts_29 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3738 = perfCnts_30 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3740 = perfCnts_31 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3742 = perfCnts_32 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3744 = perfCnts_33 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3776 = perfCnts_49 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3778 = perfCnts_50 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3780 = perfCnts_51 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3782 = perfCnts_52 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3784 = perfCnts_53 + 64'h1; // @[CSR.scala 837:71]
  wire [63:0] _T_3934 = perfCnts_2 + 64'h2; // @[CSR.scala 845:86]
  wire [64:0] _T_3935 = {{1'd0}, perfCnts_99}; // @[CSR.scala 847:69]
  wire [64:0] _T_3937 = {{1'd0}, perfCnts_100}; // @[CSR.scala 848:69]
  wire [64:0] _T_3939 = {{1'd0}, perfCnts_102}; // @[CSR.scala 849:69]
  reg [1:0] _T_4178; // @[CSR.scala 892:34]
  reg [63:0] _T_4179; // @[CSR.scala 893:34]
  reg [63:0] _T_4181; // @[CSR.scala 894:34]
  reg [63:0] _T_4182; // @[CSR.scala 895:34]
  reg [63:0] _T_4183; // @[CSR.scala 896:34]
  reg [63:0] _T_4184; // @[CSR.scala 897:34]
  reg [63:0] _T_4185; // @[CSR.scala 898:34]
  wire  _GEN_335 = _T_2885 & DISPLAY_ENABLE; // @[Debug.scala 56:24]
  wire  _GEN_337 = _T_2921 & DISPLAY_ENABLE; // @[Debug.scala 56:24]
  assign io_out_valid = io_in_valid; // @[CSR.scala 731:16]
  assign io_out_bits = _T_1490 | _T_1330; // @[CSR.scala 480:15]
  assign io_redirect_target = resetSatp ? _T_3249 : _T_3250; // @[CSR.scala 638:22]
  assign io_redirect_valid = _T_3246 | resetSatp; // @[CSR.scala 636:21]
  assign io_intrNO = raiseIntr ? causeNO : 64'h0; // @[CSR.scala 631:13]
  assign io_imemMMU_priviledgeMode = priviledgeMode; // @[CSR.scala 527:29]
  assign io_dmemMMU_priviledgeMode = mstatusStruct_mprv ? mstatusStruct_mpp : priviledgeMode; // @[CSR.scala 528:29]
  assign io_dmemMMU_status_sum = mstatus[18]; // @[CSR.scala 530:25]
  assign io_dmemMMU_status_mxr = mstatus[19]; // @[CSR.scala 532:25]
  assign io_wenFix = |raiseExceptionVec; // @[CSR.scala 628:13]
  assign _T_4181_0 = _T_4181;
  assign _T_4184_0 = _T_4184;
  assign _T_4185_0 = _T_4185;
  assign perfCnts_2_0 = perfCnts_2;
  assign satp_0 = satp;
  assign _T_4178_0 = _T_4178;
  assign intrVec_0 = intrVec;
  assign _T_4183_0 = _T_4183;
  assign _T_4182_0 = _T_4182;
  assign perfCnts_0_0 = perfCnts_0;
  assign _T_4179_0 = _T_4179;
  assign lrAddr_0 = lrAddr;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mtvec = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mcounteren = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  mcause = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  mtval = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  mepc = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  mie = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mipReg = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  misa = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  mstatus = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  medeleg = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  mideleg = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  mscratch = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  pmpcfg0 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  pmpcfg1 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  pmpcfg2 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  pmpcfg3 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  pmpaddr0 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  pmpaddr1 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  pmpaddr2 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  pmpaddr3 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  stvec = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  satp = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  sepc = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  scause = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  stval = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  sscratch = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  scounteren = _RAND_26[63:0];
  _RAND_27 = {1{`RANDOM}};
  lr = _RAND_27[0:0];
  _RAND_28 = {2{`RANDOM}};
  lrAddr = _RAND_28[63:0];
  _RAND_29 = {1{`RANDOM}};
  priviledgeMode = _RAND_29[1:0];
  _RAND_30 = {2{`RANDOM}};
  perfCnts_0 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  perfCnts_1 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  perfCnts_2 = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  perfCnts_3 = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  perfCnts_4 = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  perfCnts_5 = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  perfCnts_6 = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  perfCnts_7 = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  perfCnts_8 = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  perfCnts_9 = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  perfCnts_10 = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  perfCnts_11 = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  perfCnts_12 = _RAND_42[63:0];
  _RAND_43 = {2{`RANDOM}};
  perfCnts_13 = _RAND_43[63:0];
  _RAND_44 = {2{`RANDOM}};
  perfCnts_14 = _RAND_44[63:0];
  _RAND_45 = {2{`RANDOM}};
  perfCnts_15 = _RAND_45[63:0];
  _RAND_46 = {2{`RANDOM}};
  perfCnts_16 = _RAND_46[63:0];
  _RAND_47 = {2{`RANDOM}};
  perfCnts_17 = _RAND_47[63:0];
  _RAND_48 = {2{`RANDOM}};
  perfCnts_18 = _RAND_48[63:0];
  _RAND_49 = {2{`RANDOM}};
  perfCnts_19 = _RAND_49[63:0];
  _RAND_50 = {2{`RANDOM}};
  perfCnts_20 = _RAND_50[63:0];
  _RAND_51 = {2{`RANDOM}};
  perfCnts_21 = _RAND_51[63:0];
  _RAND_52 = {2{`RANDOM}};
  perfCnts_22 = _RAND_52[63:0];
  _RAND_53 = {2{`RANDOM}};
  perfCnts_23 = _RAND_53[63:0];
  _RAND_54 = {2{`RANDOM}};
  perfCnts_24 = _RAND_54[63:0];
  _RAND_55 = {2{`RANDOM}};
  perfCnts_25 = _RAND_55[63:0];
  _RAND_56 = {2{`RANDOM}};
  perfCnts_26 = _RAND_56[63:0];
  _RAND_57 = {2{`RANDOM}};
  perfCnts_27 = _RAND_57[63:0];
  _RAND_58 = {2{`RANDOM}};
  perfCnts_28 = _RAND_58[63:0];
  _RAND_59 = {2{`RANDOM}};
  perfCnts_29 = _RAND_59[63:0];
  _RAND_60 = {2{`RANDOM}};
  perfCnts_30 = _RAND_60[63:0];
  _RAND_61 = {2{`RANDOM}};
  perfCnts_31 = _RAND_61[63:0];
  _RAND_62 = {2{`RANDOM}};
  perfCnts_32 = _RAND_62[63:0];
  _RAND_63 = {2{`RANDOM}};
  perfCnts_33 = _RAND_63[63:0];
  _RAND_64 = {2{`RANDOM}};
  perfCnts_34 = _RAND_64[63:0];
  _RAND_65 = {2{`RANDOM}};
  perfCnts_35 = _RAND_65[63:0];
  _RAND_66 = {2{`RANDOM}};
  perfCnts_36 = _RAND_66[63:0];
  _RAND_67 = {2{`RANDOM}};
  perfCnts_37 = _RAND_67[63:0];
  _RAND_68 = {2{`RANDOM}};
  perfCnts_38 = _RAND_68[63:0];
  _RAND_69 = {2{`RANDOM}};
  perfCnts_39 = _RAND_69[63:0];
  _RAND_70 = {2{`RANDOM}};
  perfCnts_40 = _RAND_70[63:0];
  _RAND_71 = {2{`RANDOM}};
  perfCnts_41 = _RAND_71[63:0];
  _RAND_72 = {2{`RANDOM}};
  perfCnts_42 = _RAND_72[63:0];
  _RAND_73 = {2{`RANDOM}};
  perfCnts_43 = _RAND_73[63:0];
  _RAND_74 = {2{`RANDOM}};
  perfCnts_44 = _RAND_74[63:0];
  _RAND_75 = {2{`RANDOM}};
  perfCnts_45 = _RAND_75[63:0];
  _RAND_76 = {2{`RANDOM}};
  perfCnts_46 = _RAND_76[63:0];
  _RAND_77 = {2{`RANDOM}};
  perfCnts_47 = _RAND_77[63:0];
  _RAND_78 = {2{`RANDOM}};
  perfCnts_48 = _RAND_78[63:0];
  _RAND_79 = {2{`RANDOM}};
  perfCnts_49 = _RAND_79[63:0];
  _RAND_80 = {2{`RANDOM}};
  perfCnts_50 = _RAND_80[63:0];
  _RAND_81 = {2{`RANDOM}};
  perfCnts_51 = _RAND_81[63:0];
  _RAND_82 = {2{`RANDOM}};
  perfCnts_52 = _RAND_82[63:0];
  _RAND_83 = {2{`RANDOM}};
  perfCnts_53 = _RAND_83[63:0];
  _RAND_84 = {2{`RANDOM}};
  perfCnts_54 = _RAND_84[63:0];
  _RAND_85 = {2{`RANDOM}};
  perfCnts_55 = _RAND_85[63:0];
  _RAND_86 = {2{`RANDOM}};
  perfCnts_56 = _RAND_86[63:0];
  _RAND_87 = {2{`RANDOM}};
  perfCnts_57 = _RAND_87[63:0];
  _RAND_88 = {2{`RANDOM}};
  perfCnts_58 = _RAND_88[63:0];
  _RAND_89 = {2{`RANDOM}};
  perfCnts_59 = _RAND_89[63:0];
  _RAND_90 = {2{`RANDOM}};
  perfCnts_60 = _RAND_90[63:0];
  _RAND_91 = {2{`RANDOM}};
  perfCnts_61 = _RAND_91[63:0];
  _RAND_92 = {2{`RANDOM}};
  perfCnts_62 = _RAND_92[63:0];
  _RAND_93 = {2{`RANDOM}};
  perfCnts_63 = _RAND_93[63:0];
  _RAND_94 = {2{`RANDOM}};
  perfCnts_64 = _RAND_94[63:0];
  _RAND_95 = {2{`RANDOM}};
  perfCnts_65 = _RAND_95[63:0];
  _RAND_96 = {2{`RANDOM}};
  perfCnts_66 = _RAND_96[63:0];
  _RAND_97 = {2{`RANDOM}};
  perfCnts_67 = _RAND_97[63:0];
  _RAND_98 = {2{`RANDOM}};
  perfCnts_68 = _RAND_98[63:0];
  _RAND_99 = {2{`RANDOM}};
  perfCnts_69 = _RAND_99[63:0];
  _RAND_100 = {2{`RANDOM}};
  perfCnts_70 = _RAND_100[63:0];
  _RAND_101 = {2{`RANDOM}};
  perfCnts_71 = _RAND_101[63:0];
  _RAND_102 = {2{`RANDOM}};
  perfCnts_72 = _RAND_102[63:0];
  _RAND_103 = {2{`RANDOM}};
  perfCnts_73 = _RAND_103[63:0];
  _RAND_104 = {2{`RANDOM}};
  perfCnts_74 = _RAND_104[63:0];
  _RAND_105 = {2{`RANDOM}};
  perfCnts_75 = _RAND_105[63:0];
  _RAND_106 = {2{`RANDOM}};
  perfCnts_76 = _RAND_106[63:0];
  _RAND_107 = {2{`RANDOM}};
  perfCnts_77 = _RAND_107[63:0];
  _RAND_108 = {2{`RANDOM}};
  perfCnts_78 = _RAND_108[63:0];
  _RAND_109 = {2{`RANDOM}};
  perfCnts_79 = _RAND_109[63:0];
  _RAND_110 = {2{`RANDOM}};
  perfCnts_80 = _RAND_110[63:0];
  _RAND_111 = {2{`RANDOM}};
  perfCnts_81 = _RAND_111[63:0];
  _RAND_112 = {2{`RANDOM}};
  perfCnts_82 = _RAND_112[63:0];
  _RAND_113 = {2{`RANDOM}};
  perfCnts_83 = _RAND_113[63:0];
  _RAND_114 = {2{`RANDOM}};
  perfCnts_84 = _RAND_114[63:0];
  _RAND_115 = {2{`RANDOM}};
  perfCnts_85 = _RAND_115[63:0];
  _RAND_116 = {2{`RANDOM}};
  perfCnts_86 = _RAND_116[63:0];
  _RAND_117 = {2{`RANDOM}};
  perfCnts_87 = _RAND_117[63:0];
  _RAND_118 = {2{`RANDOM}};
  perfCnts_88 = _RAND_118[63:0];
  _RAND_119 = {2{`RANDOM}};
  perfCnts_89 = _RAND_119[63:0];
  _RAND_120 = {2{`RANDOM}};
  perfCnts_90 = _RAND_120[63:0];
  _RAND_121 = {2{`RANDOM}};
  perfCnts_91 = _RAND_121[63:0];
  _RAND_122 = {2{`RANDOM}};
  perfCnts_92 = _RAND_122[63:0];
  _RAND_123 = {2{`RANDOM}};
  perfCnts_93 = _RAND_123[63:0];
  _RAND_124 = {2{`RANDOM}};
  perfCnts_94 = _RAND_124[63:0];
  _RAND_125 = {2{`RANDOM}};
  perfCnts_95 = _RAND_125[63:0];
  _RAND_126 = {2{`RANDOM}};
  perfCnts_96 = _RAND_126[63:0];
  _RAND_127 = {2{`RANDOM}};
  perfCnts_97 = _RAND_127[63:0];
  _RAND_128 = {2{`RANDOM}};
  perfCnts_98 = _RAND_128[63:0];
  _RAND_129 = {2{`RANDOM}};
  perfCnts_99 = _RAND_129[63:0];
  _RAND_130 = {2{`RANDOM}};
  perfCnts_100 = _RAND_130[63:0];
  _RAND_131 = {2{`RANDOM}};
  perfCnts_101 = _RAND_131[63:0];
  _RAND_132 = {2{`RANDOM}};
  perfCnts_102 = _RAND_132[63:0];
  _RAND_133 = {2{`RANDOM}};
  perfCnts_103 = _RAND_133[63:0];
  _RAND_134 = {2{`RANDOM}};
  perfCnts_104 = _RAND_134[63:0];
  _RAND_135 = {2{`RANDOM}};
  perfCnts_105 = _RAND_135[63:0];
  _RAND_136 = {2{`RANDOM}};
  perfCnts_106 = _RAND_136[63:0];
  _RAND_137 = {2{`RANDOM}};
  perfCnts_107 = _RAND_137[63:0];
  _RAND_138 = {2{`RANDOM}};
  perfCnts_108 = _RAND_138[63:0];
  _RAND_139 = {2{`RANDOM}};
  perfCnts_109 = _RAND_139[63:0];
  _RAND_140 = {2{`RANDOM}};
  perfCnts_110 = _RAND_140[63:0];
  _RAND_141 = {2{`RANDOM}};
  perfCnts_111 = _RAND_141[63:0];
  _RAND_142 = {2{`RANDOM}};
  perfCnts_112 = _RAND_142[63:0];
  _RAND_143 = {2{`RANDOM}};
  perfCnts_113 = _RAND_143[63:0];
  _RAND_144 = {2{`RANDOM}};
  perfCnts_114 = _RAND_144[63:0];
  _RAND_145 = {2{`RANDOM}};
  perfCnts_115 = _RAND_145[63:0];
  _RAND_146 = {2{`RANDOM}};
  perfCnts_116 = _RAND_146[63:0];
  _RAND_147 = {2{`RANDOM}};
  perfCnts_117 = _RAND_147[63:0];
  _RAND_148 = {2{`RANDOM}};
  perfCnts_118 = _RAND_148[63:0];
  _RAND_149 = {2{`RANDOM}};
  perfCnts_119 = _RAND_149[63:0];
  _RAND_150 = {2{`RANDOM}};
  perfCnts_120 = _RAND_150[63:0];
  _RAND_151 = {2{`RANDOM}};
  perfCnts_121 = _RAND_151[63:0];
  _RAND_152 = {2{`RANDOM}};
  perfCnts_122 = _RAND_152[63:0];
  _RAND_153 = {2{`RANDOM}};
  perfCnts_123 = _RAND_153[63:0];
  _RAND_154 = {2{`RANDOM}};
  perfCnts_124 = _RAND_154[63:0];
  _RAND_155 = {2{`RANDOM}};
  perfCnts_125 = _RAND_155[63:0];
  _RAND_156 = {2{`RANDOM}};
  perfCnts_126 = _RAND_156[63:0];
  _RAND_157 = {2{`RANDOM}};
  perfCnts_127 = _RAND_157[63:0];
  _RAND_158 = {2{`RANDOM}};
  _T_2857 = _RAND_158[63:0];
  _RAND_159 = {2{`RANDOM}};
  _T_2866 = _RAND_159[63:0];
  _RAND_160 = {2{`RANDOM}};
  _T_2869 = _RAND_160[63:0];
  _RAND_161 = {2{`RANDOM}};
  _T_2905 = _RAND_161[63:0];
  _RAND_162 = {2{`RANDOM}};
  _T_2912 = _RAND_162[63:0];
  _RAND_163 = {2{`RANDOM}};
  _T_2926 = _RAND_163[63:0];
  _RAND_164 = {2{`RANDOM}};
  _T_2933 = _RAND_164[63:0];
  _RAND_165 = {2{`RANDOM}};
  _T_3282 = _RAND_165[63:0];
  _RAND_166 = {2{`RANDOM}};
  _T_3302 = _RAND_166[63:0];
  _RAND_167 = {2{`RANDOM}};
  _T_3311 = _RAND_167[63:0];
  _RAND_168 = {2{`RANDOM}};
  _T_3314 = _RAND_168[63:0];
  _RAND_169 = {2{`RANDOM}};
  _T_3323 = _RAND_169[63:0];
  _RAND_170 = {2{`RANDOM}};
  _T_3332 = _RAND_170[63:0];
  _RAND_171 = {1{`RANDOM}};
  _T_4178 = _RAND_171[1:0];
  _RAND_172 = {2{`RANDOM}};
  _T_4179 = _RAND_172[63:0];
  _RAND_173 = {2{`RANDOM}};
  _T_4181 = _RAND_173[63:0];
  _RAND_174 = {2{`RANDOM}};
  _T_4182 = _RAND_174[63:0];
  _RAND_175 = {2{`RANDOM}};
  _T_4183 = _RAND_175[63:0];
  _RAND_176 = {2{`RANDOM}};
  _T_4184 = _RAND_176[63:0];
  _RAND_177 = {2{`RANDOM}};
  _T_4185 = _RAND_177[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      mtvec <= 64'h0;
    end else if (_T_1908) begin
      mtvec <= wdata;
    end
    if (reset) begin
      mcounteren <= 64'h0;
    end else if (_T_1704) begin
      mcounteren <= wdata;
    end
    if (reset) begin
      mcause <= 64'h0;
    end else if (raiseExceptionIntr) begin
      if (delegS) begin
        if (_T_1680) begin
          mcause <= wdata;
        end
      end else begin
        mcause <= causeNO;
      end
    end else if (_T_1680) begin
      mcause <= wdata;
    end
    if (reset) begin
      mtval <= 64'h0;
    end else if (raiseExceptionIntr) begin
      if (delegS) begin
        if (_T_2921) begin
          mtval <= _T_2925;
        end else if (_T_2885) begin
          if (_T_2904) begin
            if (hasInstrPageFault) begin
              if (io_cfIn_crossPageIPFFix) begin
                mtval <= _T_2892;
              end else begin
                mtval <= _T_2897;
              end
            end else begin
              mtval <= _T_2902;
            end
          end else if (_T_2406) begin
            mtval <= wdata;
          end
        end else if (_T_2406) begin
          mtval <= wdata;
        end
      end else if (tvalWen) begin
        mtval <= 64'h0;
      end else if (_T_2921) begin
        mtval <= _T_2925;
      end else if (_T_2885) begin
        if (_T_2904) begin
          if (hasInstrPageFault) begin
            if (io_cfIn_crossPageIPFFix) begin
              mtval <= _T_2892;
            end else begin
              mtval <= _T_2897;
            end
          end else begin
            mtval <= _T_2902;
          end
        end else if (_T_2406) begin
          mtval <= wdata;
        end
      end else if (_T_2406) begin
        mtval <= wdata;
      end
    end else if (_T_2921) begin
      mtval <= _T_2925;
    end else if (_T_2885) begin
      if (_T_2904) begin
        if (hasInstrPageFault) begin
          if (io_cfIn_crossPageIPFFix) begin
            mtval <= _T_2892;
          end else begin
            mtval <= _T_2897;
          end
        end else begin
          mtval <= _T_2902;
        end
      end else begin
        mtval <= _GEN_144;
      end
    end else begin
      mtval <= _GEN_144;
    end
    if (raiseExceptionIntr) begin
      if (delegS) begin
        if (_T_2400) begin
          mepc <= wdata;
        end
      end else begin
        mepc <= _T_2897;
      end
    end else if (_T_2400) begin
      mepc <= wdata;
    end
    if (reset) begin
      mie <= 64'h0;
    end else if (_T_1962) begin
      mie <= wdata;
    end else if (_T_1734) begin
      mie <= _T_1738;
    end
    if (reset) begin
      mipReg <= 64'h0;
    end else if (_T_2832) begin
      mipReg <= _T_2836;
    end else if (_T_2826) begin
      mipReg <= _T_2830;
    end
    if (reset) begin
      misa <= 64'h8000000000141105;
    end else if (_T_2058) begin
      misa <= wdata;
    end
    if (reset) begin
      mstatus <= 64'h1800;
    end else if (raiseExceptionIntr) begin
      mstatus <= _T_3676;
    end else if (_T_3513) begin
      mstatus <= _T_3590;
    end else if (_T_3433) begin
      mstatus <= _T_3511;
    end else if (_T_3354) begin
      mstatus <= _T_3431;
    end else if (_T_2082) begin
      mstatus <= _T_2116;
    end else if (_T_1800) begin
      mstatus <= _T_1834;
    end
    if (reset) begin
      medeleg <= 64'h0;
    end else if (_T_1632) begin
      medeleg <= _T_1636;
    end
    if (reset) begin
      mideleg <= 64'h0;
    end else if (_T_2322) begin
      mideleg <= _T_2326;
    end
    if (reset) begin
      mscratch <= 64'h0;
    end else if (_T_2382) begin
      mscratch <= wdata;
    end
    if (reset) begin
      pmpcfg0 <= 64'h0;
    end else if (_T_2424) begin
      pmpcfg0 <= wdata;
    end
    if (reset) begin
      pmpcfg1 <= 64'h0;
    end else if (_T_2370) begin
      pmpcfg1 <= wdata;
    end
    if (reset) begin
      pmpcfg2 <= 64'h0;
    end else if (_T_1578) begin
      pmpcfg2 <= wdata;
    end
    if (reset) begin
      pmpcfg3 <= 64'h0;
    end else if (_T_2292) begin
      pmpcfg3 <= wdata;
    end
    if (reset) begin
      pmpaddr0 <= 64'h0;
    end else if (_T_2148) begin
      pmpaddr0 <= wdata;
    end
    if (reset) begin
      pmpaddr1 <= 64'h0;
    end else if (_T_1566) begin
      pmpaddr1 <= wdata;
    end
    if (reset) begin
      pmpaddr2 <= 64'h0;
    end else if (_T_2346) begin
      pmpaddr2 <= wdata;
    end
    if (reset) begin
      pmpaddr3 <= 64'h0;
    end else if (_T_1992) begin
      pmpaddr3 <= wdata;
    end
    if (reset) begin
      stvec <= 64'h0;
    end else if (_T_1650) begin
      stvec <= wdata;
    end
    if (reset) begin
      satp <= 64'h0;
    end else if (_T_1542) begin
      satp <= wdata;
    end
    if (reset) begin
      sepc <= 64'h0;
    end else if (raiseExceptionIntr) begin
      if (delegS) begin
        sepc <= _T_2897;
      end else if (_T_1668) begin
        sepc <= wdata;
      end
    end else if (_T_1668) begin
      sepc <= wdata;
    end
    if (reset) begin
      scause <= 64'h0;
    end else if (raiseExceptionIntr) begin
      if (delegS) begin
        scause <= causeNO;
      end else if (_T_2448) begin
        scause <= wdata;
      end
    end else if (_T_2448) begin
      scause <= wdata;
    end
    if (raiseExceptionIntr) begin
      if (delegS) begin
        if (tvalWen) begin
          stval <= 64'h0;
        end else if (_T_2885) begin
          if (_T_2904) begin
            if (_T_2040) begin
              stval <= wdata;
            end
          end else if (hasInstrPageFault) begin
            if (io_cfIn_crossPageIPFFix) begin
              stval <= _T_2892;
            end else begin
              stval <= _T_2897;
            end
          end else begin
            stval <= _T_2902;
          end
        end else if (_T_2040) begin
          stval <= wdata;
        end
      end else if (_T_2885) begin
        if (_T_2904) begin
          if (_T_2040) begin
            stval <= wdata;
          end
        end else begin
          stval <= _T_2903;
        end
      end else if (_T_2040) begin
        stval <= wdata;
      end
    end else if (_T_2885) begin
      if (_T_2904) begin
        stval <= _GEN_88;
      end else begin
        stval <= _T_2903;
      end
    end else begin
      stval <= _GEN_88;
    end
    if (reset) begin
      sscratch <= 64'h0;
    end else if (_T_1590) begin
      sscratch <= wdata;
    end
    if (reset) begin
      scounteren <= 64'h0;
    end else if (_T_2412) begin
      scounteren <= wdata;
    end
    if (reset) begin
      lr <= 1'h0;
    end else if (_T_3433) begin
      lr <= 1'h0;
    end else if (_T_3354) begin
      lr <= 1'h0;
    end else if (set_lr) begin
      lr <= set_lr_val;
    end
    if (reset) begin
      lrAddr <= 64'h0;
    end else if (set_lr) begin
      lrAddr <= set_lr_addr;
    end
    if (reset) begin
      priviledgeMode <= 2'h3;
    end else if (raiseExceptionIntr) begin
      if (delegS) begin
        priviledgeMode <= 2'h1;
      end else begin
        priviledgeMode <= 2'h3;
      end
    end else if (_T_3513) begin
      priviledgeMode <= 2'h0;
    end else if (_T_3433) begin
      priviledgeMode <= _T_3488;
    end else if (_T_3354) begin
      priviledgeMode <= mstatusStruct_mpp;
    end
    if (reset) begin
      perfCnts_0 <= 64'h0;
    end else begin
      perfCnts_0 <= _T_3678;
    end
    if (reset) begin
      perfCnts_1 <= 64'h0;
    end else if (_T_1968) begin
      perfCnts_1 <= wdata;
    end
    if (reset) begin
      perfCnts_2 <= 64'h0;
    end else if (perfCntCondMultiCommit) begin
      perfCnts_2 <= _T_3934;
    end else if (perfCntCondMinstret) begin
      perfCnts_2 <= _T_3682;
    end else if (_T_2286) begin
      perfCnts_2 <= wdata;
    end
    if (reset) begin
      perfCnts_3 <= 64'h0;
    end else if (perfCntCondMultiCommit) begin
      perfCnts_3 <= _T_3684;
    end else if (_T_1602) begin
      perfCnts_3 <= wdata;
    end
    if (reset) begin
      perfCnts_4 <= 64'h0;
    end else if (perfCntCondMimemStall) begin
      perfCnts_4 <= _T_3686;
    end else if (_T_1764) begin
      perfCnts_4 <= wdata;
    end
    if (reset) begin
      perfCnts_5 <= 64'h0;
    end else if (perfCntCondMaluInstr) begin
      perfCnts_5 <= _T_3688;
    end else if (_T_2190) begin
      perfCnts_5 <= wdata;
    end
    if (reset) begin
      perfCnts_6 <= 64'h0;
    end else if (perfCntCondMbruInstr) begin
      perfCnts_6 <= _T_3690;
    end else if (_T_1494) begin
      perfCnts_6 <= wdata;
    end
    if (reset) begin
      perfCnts_7 <= 64'h0;
    end else if (perfCntCondMlsuInstr) begin
      perfCnts_7 <= _T_3692;
    end else if (_T_2352) begin
      perfCnts_7 <= wdata;
    end
    if (reset) begin
      perfCnts_8 <= 64'h0;
    end else if (perfCntCondMmduInstr) begin
      perfCnts_8 <= _T_3694;
    end else if (_T_2034) begin
      perfCnts_8 <= wdata;
    end
    if (reset) begin
      perfCnts_9 <= 64'h0;
    end else if (perfCntCondMcsrInstr) begin
      perfCnts_9 <= _T_3696;
    end else if (_T_1596) begin
      perfCnts_9 <= wdata;
    end
    if (reset) begin
      perfCnts_10 <= 64'h0;
    end else if (perfCntCondMloadInstr) begin
      perfCnts_10 <= _T_3698;
    end else if (_T_1758) begin
      perfCnts_10 <= wdata;
    end
    if (reset) begin
      perfCnts_11 <= 64'h0;
    end else if (perfCntCondMmmioInstr) begin
      perfCnts_11 <= _T_3700;
    end else if (_T_1974) begin
      perfCnts_11 <= wdata;
    end
    if (reset) begin
      perfCnts_12 <= 64'h0;
    end else if (_T_2310) begin
      perfCnts_12 <= wdata;
    end
    if (reset) begin
      perfCnts_13 <= 64'h0;
    end else if (_T_1656) begin
      perfCnts_13 <= wdata;
    end
    if (reset) begin
      perfCnts_14 <= 64'h0;
    end else if (perfCntCondMmulInstr) begin
      perfCnts_14 <= _T_3706;
    end else if (_T_1842) begin
      perfCnts_14 <= wdata;
    end
    if (reset) begin
      perfCnts_15 <= 64'h0;
    end else if (perfCntCondMifuFlush) begin
      perfCnts_15 <= _T_3708;
    end else if (_T_2214) begin
      perfCnts_15 <= wdata;
    end
    if (reset) begin
      perfCnts_16 <= 64'h0;
    end else if (MbpBRight) begin
      perfCnts_16 <= _T_3710;
    end else if (_T_2478) begin
      perfCnts_16 <= wdata;
    end
    if (reset) begin
      perfCnts_17 <= 64'h0;
    end else if (MbpBWrong) begin
      perfCnts_17 <= _T_3712;
    end else if (_T_1692) begin
      perfCnts_17 <= wdata;
    end
    if (reset) begin
      perfCnts_18 <= 64'h0;
    end else if (MbpJRight) begin
      perfCnts_18 <= _T_3714;
    end else if (_T_2484) begin
      perfCnts_18 <= wdata;
    end
    if (reset) begin
      perfCnts_19 <= 64'h0;
    end else if (MbpJWrong) begin
      perfCnts_19 <= _T_3716;
    end else if (_T_2118) begin
      perfCnts_19 <= wdata;
    end
    if (reset) begin
      perfCnts_20 <= 64'h0;
    end else if (MbpIRight) begin
      perfCnts_20 <= _T_3718;
    end else if (_T_1860) begin
      perfCnts_20 <= wdata;
    end
    if (reset) begin
      perfCnts_21 <= 64'h0;
    end else if (MbpIWrong) begin
      perfCnts_21 <= _T_3720;
    end else if (_T_1530) begin
      perfCnts_21 <= wdata;
    end
    if (reset) begin
      perfCnts_22 <= 64'h0;
    end else if (MbpRRight) begin
      perfCnts_22 <= _T_3722;
    end else if (_T_2232) begin
      perfCnts_22 <= wdata;
    end
    if (reset) begin
      perfCnts_23 <= 64'h0;
    end else if (MbpRWrong) begin
      perfCnts_23 <= _T_3724;
    end else if (_T_2004) begin
      perfCnts_23 <= wdata;
    end
    if (reset) begin
      perfCnts_24 <= 64'h0;
    end else if (_T_1776) begin
      perfCnts_24 <= wdata;
    end
    if (reset) begin
      perfCnts_25 <= 64'h0;
    end else if (Custom1) begin
      perfCnts_25 <= _T_3728;
    end else if (_T_1788) begin
      perfCnts_25 <= wdata;
    end
    if (reset) begin
      perfCnts_26 <= 64'h0;
    end else if (Custom2) begin
      perfCnts_26 <= _T_3730;
    end else if (_T_2070) begin
      perfCnts_26 <= wdata;
    end
    if (reset) begin
      perfCnts_27 <= 64'h0;
    end else if (Custom3) begin
      perfCnts_27 <= _T_3732;
    end else if (_T_2238) begin
      perfCnts_27 <= wdata;
    end
    if (reset) begin
      perfCnts_28 <= 64'h0;
    end else if (Custom4) begin
      perfCnts_28 <= _T_3734;
    end else if (_T_1572) begin
      perfCnts_28 <= wdata;
    end
    if (reset) begin
      perfCnts_29 <= 64'h0;
    end else if (Custom5) begin
      perfCnts_29 <= _T_3736;
    end else if (_T_1866) begin
      perfCnts_29 <= wdata;
    end
    if (reset) begin
      perfCnts_30 <= 64'h0;
    end else if (Custom6) begin
      perfCnts_30 <= _T_3738;
    end else if (_T_2166) begin
      perfCnts_30 <= wdata;
    end
    if (reset) begin
      perfCnts_31 <= 64'h0;
    end else if (Custom7) begin
      perfCnts_31 <= _T_3740;
    end else if (_T_2430) begin
      perfCnts_31 <= wdata;
    end
    if (reset) begin
      perfCnts_32 <= 64'h0;
    end else if (Custom8) begin
      perfCnts_32 <= _T_3742;
    end else if (_T_2262) begin
      perfCnts_32 <= wdata;
    end
    if (reset) begin
      perfCnts_33 <= 64'h0;
    end else if (perfCntCondMsnnInstr) begin
      perfCnts_33 <= _T_3744;
    end else if (_T_1956) begin
      perfCnts_33 <= wdata;
    end
    if (reset) begin
      perfCnts_34 <= 64'h0;
    end else if (_T_2196) begin
      perfCnts_34 <= wdata;
    end
    if (reset) begin
      perfCnts_35 <= 64'h0;
    end else if (_T_1878) begin
      perfCnts_35 <= wdata;
    end
    if (reset) begin
      perfCnts_36 <= 64'h0;
    end else if (_T_1644) begin
      perfCnts_36 <= wdata;
    end
    if (reset) begin
      perfCnts_37 <= 64'h0;
    end else if (_T_2340) begin
      perfCnts_37 <= wdata;
    end
    if (reset) begin
      perfCnts_38 <= 64'h0;
    end else if (_T_1536) begin
      perfCnts_38 <= wdata;
    end
    if (reset) begin
      perfCnts_39 <= 64'h0;
    end else if (_T_2334) begin
      perfCnts_39 <= wdata;
    end
    if (reset) begin
      perfCnts_40 <= 64'h0;
    end else if (_T_2016) begin
      perfCnts_40 <= wdata;
    end
    if (reset) begin
      perfCnts_41 <= 64'h0;
    end else if (_T_1626) begin
      perfCnts_41 <= wdata;
    end
    if (reset) begin
      perfCnts_42 <= 64'h0;
    end else if (_T_1794) begin
      perfCnts_42 <= wdata;
    end
    if (reset) begin
      perfCnts_43 <= 64'h0;
    end else if (_T_1944) begin
      perfCnts_43 <= wdata;
    end
    if (reset) begin
      perfCnts_44 <= 64'h0;
    end else if (_T_2244) begin
      perfCnts_44 <= wdata;
    end
    if (reset) begin
      perfCnts_45 <= 64'h0;
    end else if (_T_1698) begin
      perfCnts_45 <= wdata;
    end
    if (reset) begin
      perfCnts_46 <= 64'h0;
    end else if (_T_1884) begin
      perfCnts_46 <= wdata;
    end
    if (reset) begin
      perfCnts_47 <= 64'h0;
    end else if (_T_2184) begin
      perfCnts_47 <= wdata;
    end
    if (reset) begin
      perfCnts_48 <= 64'h0;
    end else if (_T_2442) begin
      perfCnts_48 <= wdata;
    end
    if (reset) begin
      perfCnts_49 <= 64'h0;
    end else if (perfCntCondMrawStall) begin
      perfCnts_49 <= _T_3776;
    end else if (_T_2268) begin
      perfCnts_49 <= wdata;
    end
    if (reset) begin
      perfCnts_50 <= 64'h0;
    end else if (perfCntCondMexuBusy) begin
      perfCnts_50 <= _T_3778;
    end else if (_T_2472) begin
      perfCnts_50 <= wdata;
    end
    if (reset) begin
      perfCnts_51 <= 64'h0;
    end else if (perfCntCondMloadStall) begin
      perfCnts_51 <= _T_3780;
    end else if (_T_2130) begin
      perfCnts_51 <= wdata;
    end
    if (reset) begin
      perfCnts_52 <= 64'h0;
    end else if (perfCntCondMstoreStall) begin
      perfCnts_52 <= _T_3782;
    end else if (_T_1848) begin
      perfCnts_52 <= wdata;
    end
    if (reset) begin
      perfCnts_53 <= 64'h0;
    end else if (perfCntCondISUIssue) begin
      perfCnts_53 <= _T_3784;
    end else if (_T_1608) begin
      perfCnts_53 <= wdata;
    end
    if (reset) begin
      perfCnts_54 <= 64'h0;
    end else if (_T_2304) begin
      perfCnts_54 <= wdata;
    end
    if (reset) begin
      perfCnts_55 <= 64'h0;
    end else if (_T_2028) begin
      perfCnts_55 <= wdata;
    end
    if (reset) begin
      perfCnts_56 <= 64'h0;
    end else if (_T_1770) begin
      perfCnts_56 <= wdata;
    end
    if (reset) begin
      perfCnts_57 <= 64'h0;
    end else if (_T_1752) begin
      perfCnts_57 <= wdata;
    end
    if (reset) begin
      perfCnts_58 <= 64'h0;
    end else if (_T_2052) begin
      perfCnts_58 <= wdata;
    end
    if (reset) begin
      perfCnts_59 <= 64'h0;
    end else if (_T_2274) begin
      perfCnts_59 <= wdata;
    end
    if (reset) begin
      perfCnts_60 <= 64'h0;
    end else if (_T_1506) begin
      perfCnts_60 <= wdata;
    end
    if (reset) begin
      perfCnts_61 <= 64'h0;
    end else if (_T_1836) begin
      perfCnts_61 <= wdata;
    end
    if (reset) begin
      perfCnts_62 <= 64'h0;
    end else if (_T_2154) begin
      perfCnts_62 <= wdata;
    end
    if (reset) begin
      perfCnts_63 <= 64'h0;
    end else if (_T_2454) begin
      perfCnts_63 <= wdata;
    end
    if (reset) begin
      perfCnts_64 <= 64'h0;
    end else if (_T_1674) begin
      perfCnts_64 <= wdata;
    end
    if (reset) begin
      perfCnts_65 <= 64'h0;
    end else if (_T_2460) begin
      perfCnts_65 <= wdata;
    end
    if (reset) begin
      perfCnts_66 <= 64'h0;
    end else if (_T_2208) begin
      perfCnts_66 <= wdata;
    end
    if (reset) begin
      perfCnts_67 <= 64'h0;
    end else if (_T_1896) begin
      perfCnts_67 <= wdata;
    end
    if (reset) begin
      perfCnts_68 <= 64'h0;
    end else if (_T_1710) begin
      perfCnts_68 <= wdata;
    end
    if (reset) begin
      perfCnts_69 <= 64'h0;
    end else if (_T_2298) begin
      perfCnts_69 <= wdata;
    end
    if (reset) begin
      perfCnts_70 <= 64'h0;
    end else if (_T_1584) begin
      perfCnts_70 <= wdata;
    end
    if (reset) begin
      perfCnts_71 <= 64'h0;
    end else if (_T_2466) begin
      perfCnts_71 <= wdata;
    end
    if (reset) begin
      perfCnts_72 <= 64'h0;
    end else if (_T_2202) begin
      perfCnts_72 <= wdata;
    end
    if (reset) begin
      perfCnts_73 <= 64'h0;
    end else if (_T_1500) begin
      perfCnts_73 <= wdata;
    end
    if (reset) begin
      perfCnts_74 <= 64'h0;
    end else if (_T_1746) begin
      perfCnts_74 <= wdata;
    end
    if (reset) begin
      perfCnts_75 <= 64'h0;
    end else if (_T_1980) begin
      perfCnts_75 <= wdata;
    end
    if (reset) begin
      perfCnts_76 <= 64'h0;
    end else if (_T_2256) begin
      perfCnts_76 <= wdata;
    end
    if (reset) begin
      perfCnts_77 <= 64'h0;
    end else if (_T_1662) begin
      perfCnts_77 <= wdata;
    end
    if (reset) begin
      perfCnts_78 <= 64'h0;
    end else if (_T_1938) begin
      perfCnts_78 <= wdata;
    end
    if (reset) begin
      perfCnts_79 <= 64'h0;
    end else if (_T_1782) begin
      perfCnts_79 <= wdata;
    end
    if (reset) begin
      perfCnts_80 <= 64'h0;
    end else if (_T_2022) begin
      perfCnts_80 <= wdata;
    end
    if (reset) begin
      perfCnts_81 <= 64'h0;
    end else if (_T_1620) begin
      perfCnts_81 <= wdata;
    end
    if (reset) begin
      perfCnts_82 <= 64'h0;
    end else if (_T_2436) begin
      perfCnts_82 <= wdata;
    end
    if (reset) begin
      perfCnts_83 <= 64'h0;
    end else if (_T_2172) begin
      perfCnts_83 <= wdata;
    end
    if (reset) begin
      perfCnts_84 <= 64'h0;
    end else if (_T_1872) begin
      perfCnts_84 <= wdata;
    end
    if (reset) begin
      perfCnts_85 <= 64'h0;
    end else if (_T_1560) begin
      perfCnts_85 <= wdata;
    end
    if (reset) begin
      perfCnts_86 <= 64'h0;
    end else if (_T_2376) begin
      perfCnts_86 <= wdata;
    end
    if (reset) begin
      perfCnts_87 <= 64'h0;
    end else if (_T_2226) begin
      perfCnts_87 <= wdata;
    end
    if (reset) begin
      perfCnts_88 <= 64'h0;
    end else if (_T_1926) begin
      perfCnts_88 <= wdata;
    end
    if (reset) begin
      perfCnts_89 <= 64'h0;
    end else if (_T_1728) begin
      perfCnts_89 <= wdata;
    end
    if (reset) begin
      perfCnts_90 <= 64'h0;
    end else if (_T_1998) begin
      perfCnts_90 <= wdata;
    end
    if (reset) begin
      perfCnts_91 <= 64'h0;
    end else if (_T_2328) begin
      perfCnts_91 <= wdata;
    end
    if (reset) begin
      perfCnts_92 <= 64'h0;
    end else if (_T_1524) begin
      perfCnts_92 <= wdata;
    end
    if (reset) begin
      perfCnts_93 <= 64'h0;
    end else if (_T_1914) begin
      perfCnts_93 <= wdata;
    end
    if (reset) begin
      perfCnts_94 <= 64'h0;
    end else if (_T_1722) begin
      perfCnts_94 <= wdata;
    end
    if (reset) begin
      perfCnts_95 <= 64'h0;
    end else if (_T_2076) begin
      perfCnts_95 <= wdata;
    end
    if (reset) begin
      perfCnts_96 <= 64'h0;
    end else if (_T_2364) begin
      perfCnts_96 <= wdata;
    end
    if (reset) begin
      perfCnts_97 <= 64'h0;
    end else if (_T_2418) begin
      perfCnts_97 <= wdata;
    end
    if (reset) begin
      perfCnts_98 <= 64'h0;
    end else if (_T_2136) begin
      perfCnts_98 <= wdata;
    end
    if (reset) begin
      perfCnts_99 <= 64'h0;
    end else begin
      perfCnts_99 <= _T_3935[63:0];
    end
    if (reset) begin
      perfCnts_100 <= 64'h0;
    end else begin
      perfCnts_100 <= _T_3937[63:0];
    end
    if (reset) begin
      perfCnts_101 <= 64'h0;
    end else begin
      perfCnts_101 <= _T_3939[63:0];
    end
    if (reset) begin
      perfCnts_102 <= 64'h0;
    end else if (_T_1548) begin
      perfCnts_102 <= wdata;
    end
    if (reset) begin
      perfCnts_103 <= 64'h0;
    end else if (_T_2316) begin
      perfCnts_103 <= wdata;
    end
    if (reset) begin
      perfCnts_104 <= 64'h0;
    end else if (_T_2220) begin
      perfCnts_104 <= wdata;
    end
    if (reset) begin
      perfCnts_105 <= 64'h0;
    end else if (_T_1512) begin
      perfCnts_105 <= wdata;
    end
    if (reset) begin
      perfCnts_106 <= 64'h0;
    end else if (_T_1716) begin
      perfCnts_106 <= wdata;
    end
    if (reset) begin
      perfCnts_107 <= 64'h0;
    end else if (_T_2046) begin
      perfCnts_107 <= wdata;
    end
    if (reset) begin
      perfCnts_108 <= 64'h0;
    end else if (_T_2280) begin
      perfCnts_108 <= wdata;
    end
    if (reset) begin
      perfCnts_109 <= 64'h0;
    end else if (_T_1686) begin
      perfCnts_109 <= wdata;
    end
    if (reset) begin
      perfCnts_110 <= 64'h0;
    end else if (_T_1890) begin
      perfCnts_110 <= wdata;
    end
    if (reset) begin
      perfCnts_111 <= 64'h0;
    end else if (_T_2160) begin
      perfCnts_111 <= wdata;
    end
    if (reset) begin
      perfCnts_112 <= 64'h0;
    end else if (_T_2064) begin
      perfCnts_112 <= wdata;
    end
    if (reset) begin
      perfCnts_113 <= 64'h0;
    end else if (_T_1638) begin
      perfCnts_113 <= wdata;
    end
    if (reset) begin
      perfCnts_114 <= 64'h0;
    end else if (_T_2394) begin
      perfCnts_114 <= wdata;
    end
    if (reset) begin
      perfCnts_115 <= 64'h0;
    end else if (_T_2124) begin
      perfCnts_115 <= wdata;
    end
    if (reset) begin
      perfCnts_116 <= 64'h0;
    end else if (_T_1854) begin
      perfCnts_116 <= wdata;
    end
    if (reset) begin
      perfCnts_117 <= 64'h0;
    end else if (_T_1554) begin
      perfCnts_117 <= wdata;
    end
    if (reset) begin
      perfCnts_118 <= 64'h0;
    end else if (_T_2358) begin
      perfCnts_118 <= wdata;
    end
    if (reset) begin
      perfCnts_119 <= 64'h0;
    end else if (_T_1986) begin
      perfCnts_119 <= wdata;
    end
    if (reset) begin
      perfCnts_120 <= 64'h0;
    end else if (_T_1920) begin
      perfCnts_120 <= wdata;
    end
    if (reset) begin
      perfCnts_121 <= 64'h0;
    end else if (_T_1740) begin
      perfCnts_121 <= wdata;
    end
    if (reset) begin
      perfCnts_122 <= 64'h0;
    end else if (_T_1950) begin
      perfCnts_122 <= wdata;
    end
    if (reset) begin
      perfCnts_123 <= 64'h0;
    end else if (_T_2250) begin
      perfCnts_123 <= wdata;
    end
    if (reset) begin
      perfCnts_124 <= 64'h0;
    end else if (_T_1518) begin
      perfCnts_124 <= wdata;
    end
    if (reset) begin
      perfCnts_125 <= 64'h0;
    end else if (_T_1932) begin
      perfCnts_125 <= wdata;
    end
    if (reset) begin
      perfCnts_126 <= 64'h0;
    end else if (_T_2178) begin
      perfCnts_126 <= wdata;
    end
    if (reset) begin
      perfCnts_127 <= 64'h0;
    end else if (_T_2010) begin
      perfCnts_127 <= wdata;
    end
    if (reset) begin
      _T_2857 <= 64'h0;
    end else begin
      _T_2857 <= _T_2859;
    end
    if (reset) begin
      _T_2866 <= 64'h0;
    end else begin
      _T_2866 <= _T_2868;
    end
    if (reset) begin
      _T_2869 <= 64'h0;
    end else begin
      _T_2869 <= _T_2871;
    end
    if (reset) begin
      _T_2905 <= 64'h0;
    end else begin
      _T_2905 <= _T_2907;
    end
    if (reset) begin
      _T_2912 <= 64'h0;
    end else begin
      _T_2912 <= _T_2914;
    end
    if (reset) begin
      _T_2926 <= 64'h0;
    end else begin
      _T_2926 <= _T_2928;
    end
    if (reset) begin
      _T_2933 <= 64'h0;
    end else begin
      _T_2933 <= _T_2935;
    end
    if (reset) begin
      _T_3282 <= 64'h0;
    end else begin
      _T_3282 <= _T_3284;
    end
    if (reset) begin
      _T_3302 <= 64'h0;
    end else begin
      _T_3302 <= _T_3304;
    end
    if (reset) begin
      _T_3311 <= 64'h0;
    end else begin
      _T_3311 <= _T_3313;
    end
    if (reset) begin
      _T_3314 <= 64'h0;
    end else begin
      _T_3314 <= _T_3316;
    end
    if (reset) begin
      _T_3323 <= 64'h0;
    end else begin
      _T_3323 <= _T_3325;
    end
    if (reset) begin
      _T_3332 <= 64'h0;
    end else begin
      _T_3332 <= _T_3334;
    end
    _T_4178 <= priviledgeMode;
    _T_4179 <= mstatus;
    _T_4181 <= mstatus & 64'h80000003000de122;
    _T_4182 <= mepc;
    _T_4183 <= sepc;
    _T_4184 <= mcause;
    _T_4185 <= scause;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2861 & _T_2863) begin
          $fwrite(32'h80000002,"[%d] CSR: ",_T_2857); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2861 & _T_2863) begin
          $fwrite(32'h80000002,"csr write: pc %x addr %x rdata %x wdata %x func %x\n",io_cfIn_pc,addr,rdata,wdata,io_in_bits_func); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2861 & _T_2863) begin
          $fwrite(32'h80000002,"[%d] CSR: ",_T_2869); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2861 & _T_2863) begin
          $fwrite(32'h80000002,"[MST] time %d pc %x mstatus %x mideleg %x medeleg %x mode %x\n",_T_2866,io_cfIn_pc,mstatus,mideleg,medeleg,priviledgeMode); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_335 & _T_2863) begin
          $fwrite(32'h80000002,"[%d] CSR: ",_T_2912); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_335 & _T_2863) begin
          $fwrite(32'h80000002,"[PF] %d: ipf %b tval %x := addr %x pc %x priviledgeMode %x\n",_T_2905,hasInstrPageFault,_T_2903,_T_2902,io_cfIn_pc,priviledgeMode); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_337 & _T_2863) begin
          $fwrite(32'h80000002,"[%d] CSR: ",_T_2933); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_337 & _T_2863) begin
          $fwrite(32'h80000002,"[ML] %d: addr %x pc %x priviledgeMode %x\n",_T_2926,_T_2925,io_cfIn_pc,priviledgeMode); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3286 & _T_2863) begin
          $fwrite(32'h80000002,"[%d] CSR: ",_T_3282); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3286 & _T_2863) begin
          $fwrite(32'h80000002,"excin %b excgen %b",_T_3197,_T_3212); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3286 & _T_2863) begin
          $fwrite(32'h80000002,"[%d] CSR: ",_T_3302); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3286 & _T_2863) begin
          $fwrite(32'h80000002,"int/exc: pc %x int (%d):%x exc: (%d):%x\n",io_cfIn_pc,intrNO,_T_3168,exceptionNO,raiseExceptionVec); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3286 & _T_2863) begin
          $fwrite(32'h80000002,"[%d] CSR: ",_T_3314); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3286 & _T_2863) begin
          $fwrite(32'h80000002,"[MST] time %d pc %x mstatus %x mideleg %x medeleg %x mode %x\n",_T_3311,io_cfIn_pc,mstatus,mideleg,medeleg,priviledgeMode); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3327 & _T_2863) begin
          $fwrite(32'h80000002,"[%d] CSR: ",_T_3323); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3327 & _T_2863) begin
          $fwrite(32'h80000002,"redirect to %x\n",io_redirect_target); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3336 & _T_2863) begin
          $fwrite(32'h80000002,"[%d] CSR: ",_T_3332); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3336 & _T_2863) begin
          $fwrite(32'h80000002,"satp reset\n"); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"======== PerfCnt =========\n"); // @[CSR.scala 876:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- Mcycle\n",perfCnts_0); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- Minstret\n",perfCnts_2); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- MultiCommit\n",perfCnts_3); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- MimemStall\n",perfCnts_4); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- MaluInstr\n",perfCnts_5); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- MbruInstr\n",perfCnts_6); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- MlsuInstr\n",perfCnts_7); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- MmduInstr\n",perfCnts_8); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- McsrInstr\n",perfCnts_9); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- MloadInstr\n",perfCnts_10); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- MmmioInstr\n",perfCnts_11); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- MicacheHit\n",perfCnts_12); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- MdcacheHit\n",perfCnts_13); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- MmulInstr\n",perfCnts_14); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- MifuFlush\n",perfCnts_15); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- MbpBRight\n",perfCnts_16); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- MbpBWrong\n",perfCnts_17); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- MbpJRight\n",perfCnts_18); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- MbpJWrong\n",perfCnts_19); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- MbpIRight\n",perfCnts_20); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- MbpIWrong\n",perfCnts_21); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- MbpRRight\n",perfCnts_22); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- MbpRWrong\n",perfCnts_23); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- Ml2cacheHit\n",perfCnts_24); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- Custom1\n",perfCnts_25); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- Custom2\n",perfCnts_26); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- Custom3\n",perfCnts_27); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- Custom4\n",perfCnts_28); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- Custom5\n",perfCnts_29); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- Custom6\n",perfCnts_30); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- Custom7\n",perfCnts_31); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- Custom8\n",perfCnts_32); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- MsnnInstr\n",perfCnts_33); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- MrawStall\n",perfCnts_49); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- MexuBusy\n",perfCnts_50); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- MloadStall\n",perfCnts_51); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- MstoreStall\n",perfCnts_52); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d <- ISUIssue\n",perfCnts_53); // @[CSR.scala 878:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"======== PerfCntCSV =========\n\n"); // @[CSR.scala 880:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"Mcycle, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"Minstret, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"MultiCommit, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"MimemStall, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"MaluInstr, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"MbruInstr, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"MlsuInstr, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"MmduInstr, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"McsrInstr, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"MloadInstr, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"MmmioInstr, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"MicacheHit, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"MdcacheHit, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"MmulInstr, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"MifuFlush, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"MbpBRight, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"MbpBWrong, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"MbpJRight, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"MbpJWrong, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"MbpIRight, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"MbpIWrong, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"MbpRRight, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"MbpRWrong, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"Ml2cacheHit, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"Custom1, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"Custom2, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"Custom3, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"Custom4, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"Custom5, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"Custom6, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"Custom7, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"Custom8, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"MsnnInstr, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"MrawStall, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"MexuBusy, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"MloadStall, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"MstoreStall, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"ISUIssue, "); // @[CSR.scala 882:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"\n\n\n"); // @[CSR.scala 883:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_0); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_2); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_3); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_4); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_5); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_6); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_7); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_8); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_9); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_10); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_11); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_12); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_13); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_14); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_15); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_16); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_17); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_18); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_19); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_20); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_21); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_22); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_23); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_24); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_25); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_26); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_27); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_28); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_29); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_30); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_31); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_32); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_33); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_49); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_50); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_51); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_52); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"%d, ",perfCnts_53); // @[CSR.scala 885:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (nutcoretrap_0 & _T_2863) begin
          $fwrite(32'h80000002,"\n\n\n"); // @[CSR.scala 886:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module MOU(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [6:0]  io_in_bits_func,
  input  [38:0] io_cfIn_pc,
  output [38:0] io_redirect_target,
  output        io_redirect_valid,
  output        flushICache_0,
  input         DISPLAY_ENABLE,
  output        flushTLB_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  _T_2 = io_in_bits_func == 7'h1; // @[MOU.scala 52:36]
  wire  flushICache = io_in_valid & _T_2; // @[MOU.scala 52:27]
  reg [63:0] _T_3; // @[GTimer.scala 24:20]
  wire [63:0] _T_5 = _T_3 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_7 = flushICache & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  wire  _T_9 = ~reset; // @[Debug.scala 56:24]
  wire  _T_12 = io_in_bits_func == 7'h2; // @[MOU.scala 56:33]
  wire  flushTLB = io_in_valid & _T_12; // @[MOU.scala 56:24]
  reg [63:0] _T_13; // @[GTimer.scala 24:20]
  wire [63:0] _T_15 = _T_13 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_17 = flushTLB & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  assign io_redirect_target = io_cfIn_pc + 39'h4; // @[MOU.scala 49:22]
  assign io_redirect_valid = io_in_valid; // @[MOU.scala 50:21]
  assign flushICache_0 = flushICache;
  assign flushTLB_0 = flushTLB;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  _T_3 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  _T_13 = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_3 <= 64'h0;
    end else begin
      _T_3 <= _T_5;
    end
    if (reset) begin
      _T_13 <= 64'h0;
    end else begin
      _T_13 <= _T_15;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7 & _T_9) begin
          $fwrite(32'h80000002,"[%d] MOU: ",_T_3); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_7 & _T_9) begin
          $fwrite(32'h80000002,"Flush I$ at %x\n",io_cfIn_pc); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_17 & _T_9) begin
          $fwrite(32'h80000002,"[%d] MOU: ",_T_13); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_17 & _T_9) begin
          $fwrite(32'h80000002,"Sfence.vma at %x\n",io_cfIn_pc); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module SpikeProc(
  input         io_in_valid,
  input  [63:0] io_in_bits_src1,
  input  [63:0] io_in_bits_src2,
  input  [63:0] io_in_bits_op,
  output        io_out_valid,
  output [63:0] io_out_bits
);
  wire [63:0] andsRes = io_in_bits_src1 & io_in_bits_src2; // @[SpikePP.scala 37:24]
  wire [1:0] _T_64 = io_in_bits_src1[0] + io_in_bits_src1[1]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_66 = io_in_bits_src1[2] + io_in_bits_src1[3]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_68 = _T_64 + _T_66; // @[Bitwise.scala 47:55]
  wire [1:0] _T_70 = io_in_bits_src1[4] + io_in_bits_src1[5]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_72 = io_in_bits_src1[6] + io_in_bits_src1[7]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_74 = _T_70 + _T_72; // @[Bitwise.scala 47:55]
  wire [3:0] _T_76 = _T_68 + _T_74; // @[Bitwise.scala 47:55]
  wire [1:0] _T_78 = io_in_bits_src1[8] + io_in_bits_src1[9]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_80 = io_in_bits_src1[10] + io_in_bits_src1[11]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_82 = _T_78 + _T_80; // @[Bitwise.scala 47:55]
  wire [1:0] _T_84 = io_in_bits_src1[12] + io_in_bits_src1[13]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_86 = io_in_bits_src1[14] + io_in_bits_src1[15]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_88 = _T_84 + _T_86; // @[Bitwise.scala 47:55]
  wire [3:0] _T_90 = _T_82 + _T_88; // @[Bitwise.scala 47:55]
  wire [4:0] _T_92 = _T_76 + _T_90; // @[Bitwise.scala 47:55]
  wire [1:0] _T_94 = io_in_bits_src1[16] + io_in_bits_src1[17]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_96 = io_in_bits_src1[18] + io_in_bits_src1[19]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_98 = _T_94 + _T_96; // @[Bitwise.scala 47:55]
  wire [1:0] _T_100 = io_in_bits_src1[20] + io_in_bits_src1[21]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_102 = io_in_bits_src1[22] + io_in_bits_src1[23]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_104 = _T_100 + _T_102; // @[Bitwise.scala 47:55]
  wire [3:0] _T_106 = _T_98 + _T_104; // @[Bitwise.scala 47:55]
  wire [1:0] _T_108 = io_in_bits_src1[24] + io_in_bits_src1[25]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_110 = io_in_bits_src1[26] + io_in_bits_src1[27]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_112 = _T_108 + _T_110; // @[Bitwise.scala 47:55]
  wire [1:0] _T_114 = io_in_bits_src1[28] + io_in_bits_src1[29]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_116 = io_in_bits_src1[30] + io_in_bits_src1[31]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_118 = _T_114 + _T_116; // @[Bitwise.scala 47:55]
  wire [3:0] _T_120 = _T_112 + _T_118; // @[Bitwise.scala 47:55]
  wire [4:0] _T_122 = _T_106 + _T_120; // @[Bitwise.scala 47:55]
  wire [5:0] _T_124 = _T_92 + _T_122; // @[Bitwise.scala 47:55]
  wire [1:0] _T_126 = io_in_bits_src1[32] + io_in_bits_src1[33]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_128 = io_in_bits_src1[34] + io_in_bits_src1[35]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_130 = _T_126 + _T_128; // @[Bitwise.scala 47:55]
  wire [1:0] _T_132 = io_in_bits_src1[36] + io_in_bits_src1[37]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_134 = io_in_bits_src1[38] + io_in_bits_src1[39]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_136 = _T_132 + _T_134; // @[Bitwise.scala 47:55]
  wire [3:0] _T_138 = _T_130 + _T_136; // @[Bitwise.scala 47:55]
  wire [1:0] _T_140 = io_in_bits_src1[40] + io_in_bits_src1[41]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_142 = io_in_bits_src1[42] + io_in_bits_src1[43]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_144 = _T_140 + _T_142; // @[Bitwise.scala 47:55]
  wire [1:0] _T_146 = io_in_bits_src1[44] + io_in_bits_src1[45]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_148 = io_in_bits_src1[46] + io_in_bits_src1[47]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_150 = _T_146 + _T_148; // @[Bitwise.scala 47:55]
  wire [3:0] _T_152 = _T_144 + _T_150; // @[Bitwise.scala 47:55]
  wire [4:0] _T_154 = _T_138 + _T_152; // @[Bitwise.scala 47:55]
  wire [1:0] _T_156 = io_in_bits_src1[48] + io_in_bits_src1[49]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_158 = io_in_bits_src1[50] + io_in_bits_src1[51]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_160 = _T_156 + _T_158; // @[Bitwise.scala 47:55]
  wire [1:0] _T_162 = io_in_bits_src1[52] + io_in_bits_src1[53]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_164 = io_in_bits_src1[54] + io_in_bits_src1[55]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_166 = _T_162 + _T_164; // @[Bitwise.scala 47:55]
  wire [3:0] _T_168 = _T_160 + _T_166; // @[Bitwise.scala 47:55]
  wire [1:0] _T_170 = io_in_bits_src1[56] + io_in_bits_src1[57]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_172 = io_in_bits_src1[58] + io_in_bits_src1[59]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_174 = _T_170 + _T_172; // @[Bitwise.scala 47:55]
  wire [1:0] _T_176 = io_in_bits_src1[60] + io_in_bits_src1[61]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_178 = io_in_bits_src1[62] + io_in_bits_src1[63]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_180 = _T_176 + _T_178; // @[Bitwise.scala 47:55]
  wire [3:0] _T_182 = _T_174 + _T_180; // @[Bitwise.scala 47:55]
  wire [4:0] _T_184 = _T_168 + _T_182; // @[Bitwise.scala 47:55]
  wire [5:0] _T_186 = _T_154 + _T_184; // @[Bitwise.scala 47:55]
  wire [6:0] regPopRes = _T_124 + _T_186; // @[Bitwise.scala 47:55]
  wire  _T_189 = io_in_bits_op == 64'h0; // @[SpikePP.scala 36:36]
  assign io_out_valid = io_in_valid; // @[SpikePP.scala 43:18]
  assign io_out_bits = _T_189 ? andsRes : {{57'd0}, regPopRes}; // @[SpikePP.scala 40:17]
endmodule
module NeurModule(
  input         io_in_valid,
  input  [63:0] io_in_bits_src1,
  input  [63:0] io_in_bits_src2,
  input  [63:0] io_in_bits_vinit,
  input  [63:0] io_in_bits_vleak,
  input  [63:0] io_in_bits_spike,
  input  [63:0] io_in_bits_option,
  output        io_out_valid,
  output [63:0] io_out_bits
);
  wire [63:0] _GEN_0 = {{1'd0}, io_in_bits_src1[63:1]}; // @[Neuron.scala 51:27]
  wire [63:0] _T_2 = _GEN_0 + io_in_bits_src2; // @[Neuron.scala 51:27]
  wire [63:0] _T_4 = io_in_bits_vleak ^ 64'hffffffffffffffff; // @[Neuron.scala 51:55]
  wire [63:0] _T_6 = _T_4 + 64'h1; // @[Neuron.scala 51:73]
  wire [63:0] nadd = _T_2 + _T_6; // @[Neuron.scala 51:34]
  wire [64:0] naddRes = {nadd, 1'h0}; // @[Neuron.scala 52:24]
  wire  spike = _GEN_0 >= io_in_bits_src2; // @[Neuron.scala 55:29]
  wire [63:0] _T_12 = {1'h0,io_in_bits_src1[63:1]}; // @[Cat.scala 29:58]
  wire [64:0] _T_13 = {io_in_bits_src1, 1'h0}; // @[Neuron.scala 56:82]
  wire [64:0] _GEN_2 = {{64'd0}, io_in_bits_spike[0]}; // @[Neuron.scala 56:88]
  wire [64:0] _T_16 = _T_13 + _GEN_2; // @[Neuron.scala 56:88]
  wire [64:0] slsRes = io_in_bits_vinit[0] ? {{1'd0}, _T_12} : _T_16; // @[Neuron.scala 56:21]
  wire  _T_17 = io_in_bits_option == 64'h4; // @[Neuron.scala 57:38]
  wire  _T_18 = spike & _T_17; // @[Neuron.scala 57:28]
  wire  _T_19 = _T_18 & io_in_valid; // @[Neuron.scala 57:56]
  wire [63:0] _T_21 = {io_in_bits_vinit[63:1],1'h1}; // @[Cat.scala 29:58]
  wire [63:0] _T_23 = {io_in_bits_src1[63:1],1'h0}; // @[Cat.scala 29:58]
  wire [63:0] sgeRes = _T_19 ? _T_21 : _T_23; // @[Neuron.scala 57:21]
  wire  _T_24 = 64'h2 == io_in_bits_option; // @[LookupTree.scala 24:34]
  wire  _T_25 = 64'h9 == io_in_bits_option; // @[LookupTree.scala 24:34]
  wire  _T_26 = 64'h4 == io_in_bits_option; // @[LookupTree.scala 24:34]
  wire [64:0] _T_27 = _T_24 ? naddRes : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_28 = _T_25 ? slsRes : 65'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_29 = _T_26 ? sgeRes : 64'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_30 = _T_27 | _T_28; // @[Mux.scala 27:72]
  wire [64:0] _GEN_3 = {{1'd0}, _T_29}; // @[Mux.scala 27:72]
  wire [64:0] _T_31 = _T_30 | _GEN_3; // @[Mux.scala 27:72]
  assign io_out_valid = io_in_valid; // @[Neuron.scala 77:18]
  assign io_out_bits = _T_31[63:0]; // @[Neuron.scala 59:17]
endmodule
module STDP(
  input         io_in_valid,
  input  [63:0] io_in_bits_src1,
  input  [63:0] io_in_bits_src2,
  input  [63:0] io_in_bits_op,
  input  [63:0] io_in_bits_imm,
  input  [63:0] io_in_bits_output,
  input  [63:0] io_in_bits_vinit,
  output        io_out_valid,
  output [63:0] io_out_bits_res
);
  wire  stdpEnable = io_in_bits_vinit[0]; // @[STDP.scala 41:38]
  wire  _T = io_in_bits_op == 64'he; // @[STDP.scala 48:13]
  wire  _T_1 = _T & io_in_valid; // @[STDP.scala 48:33]
  wire  _T_2 = io_in_bits_op == 64'h19; // @[STDP.scala 52:19]
  wire  _T_3 = _T_2 & io_in_valid; // @[STDP.scala 52:37]
  wire  _T_4 = _T_3 & stdpEnable; // @[STDP.scala 52:46]
  wire  _T_74 = io_in_bits_src2[0] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_0 = io_in_bits_output[0] & _T_74; // @[STDP.scala 59:47]
  wire  _T_79 = io_in_bits_src2[1] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_1 = io_in_bits_output[0] & _T_79; // @[STDP.scala 59:47]
  wire  _T_84 = io_in_bits_src2[2] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_2 = io_in_bits_output[0] & _T_84; // @[STDP.scala 59:47]
  wire  _T_89 = io_in_bits_src2[3] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_3 = io_in_bits_output[0] & _T_89; // @[STDP.scala 59:47]
  wire  _T_94 = io_in_bits_src2[4] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_4 = io_in_bits_output[0] & _T_94; // @[STDP.scala 59:47]
  wire  _T_99 = io_in_bits_src2[5] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_5 = io_in_bits_output[0] & _T_99; // @[STDP.scala 59:47]
  wire  _T_104 = io_in_bits_src2[6] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_6 = io_in_bits_output[0] & _T_104; // @[STDP.scala 59:47]
  wire  _T_109 = io_in_bits_src2[7] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_7 = io_in_bits_output[0] & _T_109; // @[STDP.scala 59:47]
  wire  _T_114 = io_in_bits_src2[8] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_8 = io_in_bits_output[0] & _T_114; // @[STDP.scala 59:47]
  wire  _T_119 = io_in_bits_src2[9] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_9 = io_in_bits_output[0] & _T_119; // @[STDP.scala 59:47]
  wire  _T_124 = io_in_bits_src2[10] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_10 = io_in_bits_output[0] & _T_124; // @[STDP.scala 59:47]
  wire  _T_129 = io_in_bits_src2[11] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_11 = io_in_bits_output[0] & _T_129; // @[STDP.scala 59:47]
  wire  _T_134 = io_in_bits_src2[12] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_12 = io_in_bits_output[0] & _T_134; // @[STDP.scala 59:47]
  wire  _T_139 = io_in_bits_src2[13] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_13 = io_in_bits_output[0] & _T_139; // @[STDP.scala 59:47]
  wire  _T_144 = io_in_bits_src2[14] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_14 = io_in_bits_output[0] & _T_144; // @[STDP.scala 59:47]
  wire  _T_149 = io_in_bits_src2[15] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_15 = io_in_bits_output[0] & _T_149; // @[STDP.scala 59:47]
  wire  _T_154 = io_in_bits_src2[16] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_16 = io_in_bits_output[0] & _T_154; // @[STDP.scala 59:47]
  wire  _T_159 = io_in_bits_src2[17] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_17 = io_in_bits_output[0] & _T_159; // @[STDP.scala 59:47]
  wire  _T_164 = io_in_bits_src2[18] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_18 = io_in_bits_output[0] & _T_164; // @[STDP.scala 59:47]
  wire  _T_169 = io_in_bits_src2[19] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_19 = io_in_bits_output[0] & _T_169; // @[STDP.scala 59:47]
  wire  _T_174 = io_in_bits_src2[20] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_20 = io_in_bits_output[0] & _T_174; // @[STDP.scala 59:47]
  wire  _T_179 = io_in_bits_src2[21] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_21 = io_in_bits_output[0] & _T_179; // @[STDP.scala 59:47]
  wire  _T_184 = io_in_bits_src2[22] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_22 = io_in_bits_output[0] & _T_184; // @[STDP.scala 59:47]
  wire  _T_189 = io_in_bits_src2[23] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_23 = io_in_bits_output[0] & _T_189; // @[STDP.scala 59:47]
  wire  _T_194 = io_in_bits_src2[24] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_24 = io_in_bits_output[0] & _T_194; // @[STDP.scala 59:47]
  wire  _T_199 = io_in_bits_src2[25] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_25 = io_in_bits_output[0] & _T_199; // @[STDP.scala 59:47]
  wire  _T_204 = io_in_bits_src2[26] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_26 = io_in_bits_output[0] & _T_204; // @[STDP.scala 59:47]
  wire  _T_209 = io_in_bits_src2[27] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_27 = io_in_bits_output[0] & _T_209; // @[STDP.scala 59:47]
  wire  _T_214 = io_in_bits_src2[28] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_28 = io_in_bits_output[0] & _T_214; // @[STDP.scala 59:47]
  wire  _T_219 = io_in_bits_src2[29] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_29 = io_in_bits_output[0] & _T_219; // @[STDP.scala 59:47]
  wire  _T_224 = io_in_bits_src2[30] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_30 = io_in_bits_output[0] & _T_224; // @[STDP.scala 59:47]
  wire  _T_229 = io_in_bits_src2[31] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_31 = io_in_bits_output[0] & _T_229; // @[STDP.scala 59:47]
  wire  _T_234 = io_in_bits_src2[32] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_32 = io_in_bits_output[0] & _T_234; // @[STDP.scala 59:47]
  wire  _T_239 = io_in_bits_src2[33] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_33 = io_in_bits_output[0] & _T_239; // @[STDP.scala 59:47]
  wire  _T_244 = io_in_bits_src2[34] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_34 = io_in_bits_output[0] & _T_244; // @[STDP.scala 59:47]
  wire  _T_249 = io_in_bits_src2[35] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_35 = io_in_bits_output[0] & _T_249; // @[STDP.scala 59:47]
  wire  _T_254 = io_in_bits_src2[36] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_36 = io_in_bits_output[0] & _T_254; // @[STDP.scala 59:47]
  wire  _T_259 = io_in_bits_src2[37] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_37 = io_in_bits_output[0] & _T_259; // @[STDP.scala 59:47]
  wire  _T_264 = io_in_bits_src2[38] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_38 = io_in_bits_output[0] & _T_264; // @[STDP.scala 59:47]
  wire  _T_269 = io_in_bits_src2[39] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_39 = io_in_bits_output[0] & _T_269; // @[STDP.scala 59:47]
  wire  _T_274 = io_in_bits_src2[40] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_40 = io_in_bits_output[0] & _T_274; // @[STDP.scala 59:47]
  wire  _T_279 = io_in_bits_src2[41] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_41 = io_in_bits_output[0] & _T_279; // @[STDP.scala 59:47]
  wire  _T_284 = io_in_bits_src2[42] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_42 = io_in_bits_output[0] & _T_284; // @[STDP.scala 59:47]
  wire  _T_289 = io_in_bits_src2[43] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_43 = io_in_bits_output[0] & _T_289; // @[STDP.scala 59:47]
  wire  _T_294 = io_in_bits_src2[44] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_44 = io_in_bits_output[0] & _T_294; // @[STDP.scala 59:47]
  wire  _T_299 = io_in_bits_src2[45] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_45 = io_in_bits_output[0] & _T_299; // @[STDP.scala 59:47]
  wire  _T_304 = io_in_bits_src2[46] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_46 = io_in_bits_output[0] & _T_304; // @[STDP.scala 59:47]
  wire  _T_309 = io_in_bits_src2[47] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_47 = io_in_bits_output[0] & _T_309; // @[STDP.scala 59:47]
  wire  _T_314 = io_in_bits_src2[48] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_48 = io_in_bits_output[0] & _T_314; // @[STDP.scala 59:47]
  wire  _T_319 = io_in_bits_src2[49] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_49 = io_in_bits_output[0] & _T_319; // @[STDP.scala 59:47]
  wire  _T_324 = io_in_bits_src2[50] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_50 = io_in_bits_output[0] & _T_324; // @[STDP.scala 59:47]
  wire  _T_329 = io_in_bits_src2[51] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_51 = io_in_bits_output[0] & _T_329; // @[STDP.scala 59:47]
  wire  _T_334 = io_in_bits_src2[52] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_52 = io_in_bits_output[0] & _T_334; // @[STDP.scala 59:47]
  wire  _T_339 = io_in_bits_src2[53] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_53 = io_in_bits_output[0] & _T_339; // @[STDP.scala 59:47]
  wire  _T_344 = io_in_bits_src2[54] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_54 = io_in_bits_output[0] & _T_344; // @[STDP.scala 59:47]
  wire  _T_349 = io_in_bits_src2[55] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_55 = io_in_bits_output[0] & _T_349; // @[STDP.scala 59:47]
  wire  _T_354 = io_in_bits_src2[56] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_56 = io_in_bits_output[0] & _T_354; // @[STDP.scala 59:47]
  wire  _T_359 = io_in_bits_src2[57] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_57 = io_in_bits_output[0] & _T_359; // @[STDP.scala 59:47]
  wire  _T_364 = io_in_bits_src2[58] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_58 = io_in_bits_output[0] & _T_364; // @[STDP.scala 59:47]
  wire  _T_369 = io_in_bits_src2[59] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_59 = io_in_bits_output[0] & _T_369; // @[STDP.scala 59:47]
  wire  _T_374 = io_in_bits_src2[60] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_60 = io_in_bits_output[0] & _T_374; // @[STDP.scala 59:47]
  wire  _T_379 = io_in_bits_src2[61] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_61 = io_in_bits_output[0] & _T_379; // @[STDP.scala 59:47]
  wire  _T_384 = io_in_bits_src2[62] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_62 = io_in_bits_output[0] & _T_384; // @[STDP.scala 59:47]
  wire  _T_389 = io_in_bits_src2[63] & io_in_bits_output[0]; // @[STDP.scala 60:43]
  wire  _GEN_63 = io_in_bits_output[0] & _T_389; // @[STDP.scala 59:47]
  wire [7:0] _T_396 = {_GEN_7,_GEN_6,_GEN_5,_GEN_4,_GEN_3,_GEN_2,_GEN_1,_GEN_0}; // @[STDP.scala 63:36]
  wire [15:0] _T_404 = {_GEN_15,_GEN_14,_GEN_13,_GEN_12,_GEN_11,_GEN_10,_GEN_9,_GEN_8,_T_396}; // @[STDP.scala 63:36]
  wire [7:0] _T_411 = {_GEN_23,_GEN_22,_GEN_21,_GEN_20,_GEN_19,_GEN_18,_GEN_17,_GEN_16}; // @[STDP.scala 63:36]
  wire [31:0] _T_420 = {_GEN_31,_GEN_30,_GEN_29,_GEN_28,_GEN_27,_GEN_26,_GEN_25,_GEN_24,_T_411,_T_404}; // @[STDP.scala 63:36]
  wire [7:0] _T_427 = {_GEN_39,_GEN_38,_GEN_37,_GEN_36,_GEN_35,_GEN_34,_GEN_33,_GEN_32}; // @[STDP.scala 63:36]
  wire [15:0] _T_435 = {_GEN_47,_GEN_46,_GEN_45,_GEN_44,_GEN_43,_GEN_42,_GEN_41,_GEN_40,_T_427}; // @[STDP.scala 63:36]
  wire [7:0] _T_442 = {_GEN_55,_GEN_54,_GEN_53,_GEN_52,_GEN_51,_GEN_50,_GEN_49,_GEN_48}; // @[STDP.scala 63:36]
  wire [31:0] _T_451 = {_GEN_63,_GEN_62,_GEN_61,_GEN_60,_GEN_59,_GEN_58,_GEN_57,_GEN_56,_T_442,_T_435}; // @[STDP.scala 63:36]
  wire [63:0] _T_452 = {_T_451,_T_420}; // @[STDP.scala 63:36]
  wire [63:0] _GEN_70 = _T_4 ? _T_452 : io_in_bits_src1; // @[STDP.scala 52:60]
  assign io_out_valid = io_in_valid; // @[STDP.scala 51:22 STDP.scala 65:22 STDP.scala 69:22 STDP.scala 73:22]
  assign io_out_bits_res = _T_1 ? io_in_bits_imm : _GEN_70; // @[STDP.scala 49:25 STDP.scala 63:25 STDP.scala 67:25 STDP.scala 71:25]
endmodule
module MaxPeriodFibonacciLFSR(
  input   clock,
  input   reset,
  output  io_out_0,
  output  io_out_1,
  output  io_out_2,
  output  io_out_3,
  output  io_out_4,
  output  io_out_5,
  output  io_out_6,
  output  io_out_7,
  output  io_out_8,
  output  io_out_9,
  output  io_out_10,
  output  io_out_11,
  output  io_out_12,
  output  io_out_13,
  output  io_out_14,
  output  io_out_15
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg  state_0; // @[PRNG.scala 47:50]
  reg  state_1; // @[PRNG.scala 47:50]
  reg  state_2; // @[PRNG.scala 47:50]
  reg  state_3; // @[PRNG.scala 47:50]
  reg  state_4; // @[PRNG.scala 47:50]
  reg  state_5; // @[PRNG.scala 47:50]
  reg  state_6; // @[PRNG.scala 47:50]
  reg  state_7; // @[PRNG.scala 47:50]
  reg  state_8; // @[PRNG.scala 47:50]
  reg  state_9; // @[PRNG.scala 47:50]
  reg  state_10; // @[PRNG.scala 47:50]
  reg  state_11; // @[PRNG.scala 47:50]
  reg  state_12; // @[PRNG.scala 47:50]
  reg  state_13; // @[PRNG.scala 47:50]
  reg  state_14; // @[PRNG.scala 47:50]
  reg  state_15; // @[PRNG.scala 47:50]
  wire  _T_1 = state_15 ^ state_13; // @[LFSR.scala 15:41]
  wire  _T_2 = _T_1 ^ state_12; // @[LFSR.scala 15:41]
  wire  _T_3 = _T_2 ^ state_10; // @[LFSR.scala 15:41]
  assign io_out_0 = state_0; // @[PRNG.scala 69:10]
  assign io_out_1 = state_1; // @[PRNG.scala 69:10]
  assign io_out_2 = state_2; // @[PRNG.scala 69:10]
  assign io_out_3 = state_3; // @[PRNG.scala 69:10]
  assign io_out_4 = state_4; // @[PRNG.scala 69:10]
  assign io_out_5 = state_5; // @[PRNG.scala 69:10]
  assign io_out_6 = state_6; // @[PRNG.scala 69:10]
  assign io_out_7 = state_7; // @[PRNG.scala 69:10]
  assign io_out_8 = state_8; // @[PRNG.scala 69:10]
  assign io_out_9 = state_9; // @[PRNG.scala 69:10]
  assign io_out_10 = state_10; // @[PRNG.scala 69:10]
  assign io_out_11 = state_11; // @[PRNG.scala 69:10]
  assign io_out_12 = state_12; // @[PRNG.scala 69:10]
  assign io_out_13 = state_13; // @[PRNG.scala 69:10]
  assign io_out_14 = state_14; // @[PRNG.scala 69:10]
  assign io_out_15 = state_15; // @[PRNG.scala 69:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  state_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  state_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  state_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  state_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  state_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  state_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  state_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  state_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  state_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  state_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  state_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  state_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  state_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  state_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  state_15 = _RAND_15[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state_0 <= 1'h0;
    end else begin
      state_0 <= _T_3;
    end
    if (reset) begin
      state_1 <= 1'h0;
    end else begin
      state_1 <= state_0;
    end
    if (reset) begin
      state_2 <= 1'h0;
    end else begin
      state_2 <= state_1;
    end
    if (reset) begin
      state_3 <= 1'h0;
    end else begin
      state_3 <= state_2;
    end
    if (reset) begin
      state_4 <= 1'h0;
    end else begin
      state_4 <= state_3;
    end
    if (reset) begin
      state_5 <= 1'h0;
    end else begin
      state_5 <= state_4;
    end
    if (reset) begin
      state_6 <= 1'h0;
    end else begin
      state_6 <= state_5;
    end
    if (reset) begin
      state_7 <= 1'h0;
    end else begin
      state_7 <= state_6;
    end
    if (reset) begin
      state_8 <= 1'h0;
    end else begin
      state_8 <= state_7;
    end
    if (reset) begin
      state_9 <= 1'h0;
    end else begin
      state_9 <= state_8;
    end
    if (reset) begin
      state_10 <= 1'h0;
    end else begin
      state_10 <= state_9;
    end
    if (reset) begin
      state_11 <= 1'h0;
    end else begin
      state_11 <= state_10;
    end
    if (reset) begin
      state_12 <= 1'h0;
    end else begin
      state_12 <= state_11;
    end
    if (reset) begin
      state_13 <= 1'h0;
    end else begin
      state_13 <= state_12;
    end
    if (reset) begin
      state_14 <= 1'h0;
    end else begin
      state_14 <= state_13;
    end
    state_15 <= reset | state_14;
  end
endmodule
module LTD(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [63:0] io_in_bits_prob,
  input  [63:0] io_in_bits_syn,
  output        io_out_valid,
  output [63:0] io_out_bits_res,
  output [63:0] io_out_bits_ret,
  output [63:0] io_out_bits_cnt
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  MaxPeriodFibonacciLFSR_clock; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_reset; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_0; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_1; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_2; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_3; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_4; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_5; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_6; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_7; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_8; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_9; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_10; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_11; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_12; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_13; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_14; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_15; // @[PRNG.scala 82:22]
  reg [63:0] syn; // @[LTD.scala 40:22]
  reg [9:0] r; // @[LTD.scala 43:20]
  reg [5:0] value; // @[Counter.scala 29:33]
  reg [1:0] state; // @[LTD.scala 49:24]
  wire  _T_64 = state == 2'h0; // @[LTD.scala 50:23]
  wire  _T_65 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire  busy = _T_64 & _T_65; // @[LTD.scala 50:35]
  wire  _T_67 = state == 2'h1; // @[LTD.scala 55:22]
  wire [7:0] _T_74 = {MaxPeriodFibonacciLFSR_io_out_7,MaxPeriodFibonacciLFSR_io_out_6,MaxPeriodFibonacciLFSR_io_out_5,MaxPeriodFibonacciLFSR_io_out_4,MaxPeriodFibonacciLFSR_io_out_3,MaxPeriodFibonacciLFSR_io_out_2,MaxPeriodFibonacciLFSR_io_out_1,MaxPeriodFibonacciLFSR_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] _T_82 = {MaxPeriodFibonacciLFSR_io_out_15,MaxPeriodFibonacciLFSR_io_out_14,MaxPeriodFibonacciLFSR_io_out_13,MaxPeriodFibonacciLFSR_io_out_12,MaxPeriodFibonacciLFSR_io_out_11,MaxPeriodFibonacciLFSR_io_out_10,MaxPeriodFibonacciLFSR_io_out_9,MaxPeriodFibonacciLFSR_io_out_8,_T_74}; // @[PRNG.scala 86:17]
  wire [7:0] _T_106 = {_T_82[8],_T_82[9],_T_82[10],_T_82[11],_T_82[12],_T_82[13],_T_82[14],_T_82[15]}; // @[LFSR.scala 43:8]
  wire [15:0] _T_114 = {_T_82[0],_T_82[1],_T_82[2],_T_82[3],_T_82[4],_T_82[5],_T_82[6],_T_82[7],_T_106}; // @[LFSR.scala 43:8]
  wire [9:0] _T_117 = {_T_114[14:10],_T_114[7:3]}; // @[Cat.scala 29:58]
  wire  _T_118 = state == 2'h2; // @[LTD.scala 59:22]
  wire [63:0] _T_119 = syn >> value; // @[LTD.scala 60:17]
  wire [63:0] _GEN_340 = {{54'd0}, r}; // @[LTD.scala 61:37]
  wire  _T_122 = _GEN_340 >= io_in_bits_prob; // @[LTD.scala 61:37]
  wire  _GEN_1 = 6'h0 == value ? _T_122 : syn[0]; // @[LTD.scala 61:32]
  wire  _GEN_2 = 6'h1 == value ? _T_122 : syn[1]; // @[LTD.scala 61:32]
  wire  _GEN_3 = 6'h2 == value ? _T_122 : syn[2]; // @[LTD.scala 61:32]
  wire  _GEN_4 = 6'h3 == value ? _T_122 : syn[3]; // @[LTD.scala 61:32]
  wire  _GEN_5 = 6'h4 == value ? _T_122 : syn[4]; // @[LTD.scala 61:32]
  wire  _GEN_6 = 6'h5 == value ? _T_122 : syn[5]; // @[LTD.scala 61:32]
  wire  _GEN_7 = 6'h6 == value ? _T_122 : syn[6]; // @[LTD.scala 61:32]
  wire  _GEN_8 = 6'h7 == value ? _T_122 : syn[7]; // @[LTD.scala 61:32]
  wire  _GEN_9 = 6'h8 == value ? _T_122 : syn[8]; // @[LTD.scala 61:32]
  wire  _GEN_10 = 6'h9 == value ? _T_122 : syn[9]; // @[LTD.scala 61:32]
  wire  _GEN_11 = 6'ha == value ? _T_122 : syn[10]; // @[LTD.scala 61:32]
  wire  _GEN_12 = 6'hb == value ? _T_122 : syn[11]; // @[LTD.scala 61:32]
  wire  _GEN_13 = 6'hc == value ? _T_122 : syn[12]; // @[LTD.scala 61:32]
  wire  _GEN_14 = 6'hd == value ? _T_122 : syn[13]; // @[LTD.scala 61:32]
  wire  _GEN_15 = 6'he == value ? _T_122 : syn[14]; // @[LTD.scala 61:32]
  wire  _GEN_16 = 6'hf == value ? _T_122 : syn[15]; // @[LTD.scala 61:32]
  wire  _GEN_17 = 6'h10 == value ? _T_122 : syn[16]; // @[LTD.scala 61:32]
  wire  _GEN_18 = 6'h11 == value ? _T_122 : syn[17]; // @[LTD.scala 61:32]
  wire  _GEN_19 = 6'h12 == value ? _T_122 : syn[18]; // @[LTD.scala 61:32]
  wire  _GEN_20 = 6'h13 == value ? _T_122 : syn[19]; // @[LTD.scala 61:32]
  wire  _GEN_21 = 6'h14 == value ? _T_122 : syn[20]; // @[LTD.scala 61:32]
  wire  _GEN_22 = 6'h15 == value ? _T_122 : syn[21]; // @[LTD.scala 61:32]
  wire  _GEN_23 = 6'h16 == value ? _T_122 : syn[22]; // @[LTD.scala 61:32]
  wire  _GEN_24 = 6'h17 == value ? _T_122 : syn[23]; // @[LTD.scala 61:32]
  wire  _GEN_25 = 6'h18 == value ? _T_122 : syn[24]; // @[LTD.scala 61:32]
  wire  _GEN_26 = 6'h19 == value ? _T_122 : syn[25]; // @[LTD.scala 61:32]
  wire  _GEN_27 = 6'h1a == value ? _T_122 : syn[26]; // @[LTD.scala 61:32]
  wire  _GEN_28 = 6'h1b == value ? _T_122 : syn[27]; // @[LTD.scala 61:32]
  wire  _GEN_29 = 6'h1c == value ? _T_122 : syn[28]; // @[LTD.scala 61:32]
  wire  _GEN_30 = 6'h1d == value ? _T_122 : syn[29]; // @[LTD.scala 61:32]
  wire  _GEN_31 = 6'h1e == value ? _T_122 : syn[30]; // @[LTD.scala 61:32]
  wire  _GEN_32 = 6'h1f == value ? _T_122 : syn[31]; // @[LTD.scala 61:32]
  wire  _GEN_33 = 6'h20 == value ? _T_122 : syn[32]; // @[LTD.scala 61:32]
  wire  _GEN_34 = 6'h21 == value ? _T_122 : syn[33]; // @[LTD.scala 61:32]
  wire  _GEN_35 = 6'h22 == value ? _T_122 : syn[34]; // @[LTD.scala 61:32]
  wire  _GEN_36 = 6'h23 == value ? _T_122 : syn[35]; // @[LTD.scala 61:32]
  wire  _GEN_37 = 6'h24 == value ? _T_122 : syn[36]; // @[LTD.scala 61:32]
  wire  _GEN_38 = 6'h25 == value ? _T_122 : syn[37]; // @[LTD.scala 61:32]
  wire  _GEN_39 = 6'h26 == value ? _T_122 : syn[38]; // @[LTD.scala 61:32]
  wire  _GEN_40 = 6'h27 == value ? _T_122 : syn[39]; // @[LTD.scala 61:32]
  wire  _GEN_41 = 6'h28 == value ? _T_122 : syn[40]; // @[LTD.scala 61:32]
  wire  _GEN_42 = 6'h29 == value ? _T_122 : syn[41]; // @[LTD.scala 61:32]
  wire  _GEN_43 = 6'h2a == value ? _T_122 : syn[42]; // @[LTD.scala 61:32]
  wire  _GEN_44 = 6'h2b == value ? _T_122 : syn[43]; // @[LTD.scala 61:32]
  wire  _GEN_45 = 6'h2c == value ? _T_122 : syn[44]; // @[LTD.scala 61:32]
  wire  _GEN_46 = 6'h2d == value ? _T_122 : syn[45]; // @[LTD.scala 61:32]
  wire  _GEN_47 = 6'h2e == value ? _T_122 : syn[46]; // @[LTD.scala 61:32]
  wire  _GEN_48 = 6'h2f == value ? _T_122 : syn[47]; // @[LTD.scala 61:32]
  wire  _GEN_49 = 6'h30 == value ? _T_122 : syn[48]; // @[LTD.scala 61:32]
  wire  _GEN_50 = 6'h31 == value ? _T_122 : syn[49]; // @[LTD.scala 61:32]
  wire  _GEN_51 = 6'h32 == value ? _T_122 : syn[50]; // @[LTD.scala 61:32]
  wire  _GEN_52 = 6'h33 == value ? _T_122 : syn[51]; // @[LTD.scala 61:32]
  wire  _GEN_53 = 6'h34 == value ? _T_122 : syn[52]; // @[LTD.scala 61:32]
  wire  _GEN_54 = 6'h35 == value ? _T_122 : syn[53]; // @[LTD.scala 61:32]
  wire  _GEN_55 = 6'h36 == value ? _T_122 : syn[54]; // @[LTD.scala 61:32]
  wire  _GEN_56 = 6'h37 == value ? _T_122 : syn[55]; // @[LTD.scala 61:32]
  wire  _GEN_57 = 6'h38 == value ? _T_122 : syn[56]; // @[LTD.scala 61:32]
  wire  _GEN_58 = 6'h39 == value ? _T_122 : syn[57]; // @[LTD.scala 61:32]
  wire  _GEN_59 = 6'h3a == value ? _T_122 : syn[58]; // @[LTD.scala 61:32]
  wire  _GEN_60 = 6'h3b == value ? _T_122 : syn[59]; // @[LTD.scala 61:32]
  wire  _GEN_61 = 6'h3c == value ? _T_122 : syn[60]; // @[LTD.scala 61:32]
  wire  _GEN_62 = 6'h3d == value ? _T_122 : syn[61]; // @[LTD.scala 61:32]
  wire  _GEN_63 = 6'h3e == value ? _T_122 : syn[62]; // @[LTD.scala 61:32]
  wire  _GEN_64 = 6'h3f == value ? _T_122 : syn[63]; // @[LTD.scala 61:32]
  wire  _GEN_65 = _T_119[0] ? _GEN_1 : syn[0]; // @[LTD.scala 60:37]
  wire  _GEN_66 = _T_119[0] ? _GEN_2 : syn[1]; // @[LTD.scala 60:37]
  wire  _GEN_67 = _T_119[0] ? _GEN_3 : syn[2]; // @[LTD.scala 60:37]
  wire  _GEN_68 = _T_119[0] ? _GEN_4 : syn[3]; // @[LTD.scala 60:37]
  wire  _GEN_69 = _T_119[0] ? _GEN_5 : syn[4]; // @[LTD.scala 60:37]
  wire  _GEN_70 = _T_119[0] ? _GEN_6 : syn[5]; // @[LTD.scala 60:37]
  wire  _GEN_71 = _T_119[0] ? _GEN_7 : syn[6]; // @[LTD.scala 60:37]
  wire  _GEN_72 = _T_119[0] ? _GEN_8 : syn[7]; // @[LTD.scala 60:37]
  wire  _GEN_73 = _T_119[0] ? _GEN_9 : syn[8]; // @[LTD.scala 60:37]
  wire  _GEN_74 = _T_119[0] ? _GEN_10 : syn[9]; // @[LTD.scala 60:37]
  wire  _GEN_75 = _T_119[0] ? _GEN_11 : syn[10]; // @[LTD.scala 60:37]
  wire  _GEN_76 = _T_119[0] ? _GEN_12 : syn[11]; // @[LTD.scala 60:37]
  wire  _GEN_77 = _T_119[0] ? _GEN_13 : syn[12]; // @[LTD.scala 60:37]
  wire  _GEN_78 = _T_119[0] ? _GEN_14 : syn[13]; // @[LTD.scala 60:37]
  wire  _GEN_79 = _T_119[0] ? _GEN_15 : syn[14]; // @[LTD.scala 60:37]
  wire  _GEN_80 = _T_119[0] ? _GEN_16 : syn[15]; // @[LTD.scala 60:37]
  wire  _GEN_81 = _T_119[0] ? _GEN_17 : syn[16]; // @[LTD.scala 60:37]
  wire  _GEN_82 = _T_119[0] ? _GEN_18 : syn[17]; // @[LTD.scala 60:37]
  wire  _GEN_83 = _T_119[0] ? _GEN_19 : syn[18]; // @[LTD.scala 60:37]
  wire  _GEN_84 = _T_119[0] ? _GEN_20 : syn[19]; // @[LTD.scala 60:37]
  wire  _GEN_85 = _T_119[0] ? _GEN_21 : syn[20]; // @[LTD.scala 60:37]
  wire  _GEN_86 = _T_119[0] ? _GEN_22 : syn[21]; // @[LTD.scala 60:37]
  wire  _GEN_87 = _T_119[0] ? _GEN_23 : syn[22]; // @[LTD.scala 60:37]
  wire  _GEN_88 = _T_119[0] ? _GEN_24 : syn[23]; // @[LTD.scala 60:37]
  wire  _GEN_89 = _T_119[0] ? _GEN_25 : syn[24]; // @[LTD.scala 60:37]
  wire  _GEN_90 = _T_119[0] ? _GEN_26 : syn[25]; // @[LTD.scala 60:37]
  wire  _GEN_91 = _T_119[0] ? _GEN_27 : syn[26]; // @[LTD.scala 60:37]
  wire  _GEN_92 = _T_119[0] ? _GEN_28 : syn[27]; // @[LTD.scala 60:37]
  wire  _GEN_93 = _T_119[0] ? _GEN_29 : syn[28]; // @[LTD.scala 60:37]
  wire  _GEN_94 = _T_119[0] ? _GEN_30 : syn[29]; // @[LTD.scala 60:37]
  wire  _GEN_95 = _T_119[0] ? _GEN_31 : syn[30]; // @[LTD.scala 60:37]
  wire  _GEN_96 = _T_119[0] ? _GEN_32 : syn[31]; // @[LTD.scala 60:37]
  wire  _GEN_97 = _T_119[0] ? _GEN_33 : syn[32]; // @[LTD.scala 60:37]
  wire  _GEN_98 = _T_119[0] ? _GEN_34 : syn[33]; // @[LTD.scala 60:37]
  wire  _GEN_99 = _T_119[0] ? _GEN_35 : syn[34]; // @[LTD.scala 60:37]
  wire  _GEN_100 = _T_119[0] ? _GEN_36 : syn[35]; // @[LTD.scala 60:37]
  wire  _GEN_101 = _T_119[0] ? _GEN_37 : syn[36]; // @[LTD.scala 60:37]
  wire  _GEN_102 = _T_119[0] ? _GEN_38 : syn[37]; // @[LTD.scala 60:37]
  wire  _GEN_103 = _T_119[0] ? _GEN_39 : syn[38]; // @[LTD.scala 60:37]
  wire  _GEN_104 = _T_119[0] ? _GEN_40 : syn[39]; // @[LTD.scala 60:37]
  wire  _GEN_105 = _T_119[0] ? _GEN_41 : syn[40]; // @[LTD.scala 60:37]
  wire  _GEN_106 = _T_119[0] ? _GEN_42 : syn[41]; // @[LTD.scala 60:37]
  wire  _GEN_107 = _T_119[0] ? _GEN_43 : syn[42]; // @[LTD.scala 60:37]
  wire  _GEN_108 = _T_119[0] ? _GEN_44 : syn[43]; // @[LTD.scala 60:37]
  wire  _GEN_109 = _T_119[0] ? _GEN_45 : syn[44]; // @[LTD.scala 60:37]
  wire  _GEN_110 = _T_119[0] ? _GEN_46 : syn[45]; // @[LTD.scala 60:37]
  wire  _GEN_111 = _T_119[0] ? _GEN_47 : syn[46]; // @[LTD.scala 60:37]
  wire  _GEN_112 = _T_119[0] ? _GEN_48 : syn[47]; // @[LTD.scala 60:37]
  wire  _GEN_113 = _T_119[0] ? _GEN_49 : syn[48]; // @[LTD.scala 60:37]
  wire  _GEN_114 = _T_119[0] ? _GEN_50 : syn[49]; // @[LTD.scala 60:37]
  wire  _GEN_115 = _T_119[0] ? _GEN_51 : syn[50]; // @[LTD.scala 60:37]
  wire  _GEN_116 = _T_119[0] ? _GEN_52 : syn[51]; // @[LTD.scala 60:37]
  wire  _GEN_117 = _T_119[0] ? _GEN_53 : syn[52]; // @[LTD.scala 60:37]
  wire  _GEN_118 = _T_119[0] ? _GEN_54 : syn[53]; // @[LTD.scala 60:37]
  wire  _GEN_119 = _T_119[0] ? _GEN_55 : syn[54]; // @[LTD.scala 60:37]
  wire  _GEN_120 = _T_119[0] ? _GEN_56 : syn[55]; // @[LTD.scala 60:37]
  wire  _GEN_121 = _T_119[0] ? _GEN_57 : syn[56]; // @[LTD.scala 60:37]
  wire  _GEN_122 = _T_119[0] ? _GEN_58 : syn[57]; // @[LTD.scala 60:37]
  wire  _GEN_123 = _T_119[0] ? _GEN_59 : syn[58]; // @[LTD.scala 60:37]
  wire  _GEN_124 = _T_119[0] ? _GEN_60 : syn[59]; // @[LTD.scala 60:37]
  wire  _GEN_125 = _T_119[0] ? _GEN_61 : syn[60]; // @[LTD.scala 60:37]
  wire  _GEN_126 = _T_119[0] ? _GEN_62 : syn[61]; // @[LTD.scala 60:37]
  wire  _GEN_127 = _T_119[0] ? _GEN_63 : syn[62]; // @[LTD.scala 60:37]
  wire  _GEN_128 = _T_119[0] ? _GEN_64 : syn[63]; // @[LTD.scala 60:37]
  wire  _T_123 = value == 6'h3f; // @[Counter.scala 38:24]
  wire [5:0] _T_125 = value + 6'h1; // @[Counter.scala 39:22]
  wire  _T_126 = value != 6'h3f; // @[LTD.scala 64:24]
  wire  _GEN_135 = _T_118 ? _GEN_66 : syn[1]; // @[LTD.scala 59:33]
  wire  _GEN_205 = _T_67 ? syn[1] : _GEN_135; // @[LTD.scala 55:33]
  wire  syn_new_1 = busy ? syn[1] : _GEN_205; // @[LTD.scala 52:15]
  wire  _GEN_134 = _T_118 ? _GEN_65 : syn[0]; // @[LTD.scala 59:33]
  wire  _GEN_204 = _T_67 ? syn[0] : _GEN_134; // @[LTD.scala 55:33]
  wire  syn_new_0 = busy ? syn[0] : _GEN_204; // @[LTD.scala 52:15]
  wire  _GEN_137 = _T_118 ? _GEN_68 : syn[3]; // @[LTD.scala 59:33]
  wire  _GEN_207 = _T_67 ? syn[3] : _GEN_137; // @[LTD.scala 55:33]
  wire  syn_new_3 = busy ? syn[3] : _GEN_207; // @[LTD.scala 52:15]
  wire  _GEN_136 = _T_118 ? _GEN_67 : syn[2]; // @[LTD.scala 59:33]
  wire  _GEN_206 = _T_67 ? syn[2] : _GEN_136; // @[LTD.scala 55:33]
  wire  syn_new_2 = busy ? syn[2] : _GEN_206; // @[LTD.scala 52:15]
  wire  _GEN_139 = _T_118 ? _GEN_70 : syn[5]; // @[LTD.scala 59:33]
  wire  _GEN_209 = _T_67 ? syn[5] : _GEN_139; // @[LTD.scala 55:33]
  wire  syn_new_5 = busy ? syn[5] : _GEN_209; // @[LTD.scala 52:15]
  wire  _GEN_138 = _T_118 ? _GEN_69 : syn[4]; // @[LTD.scala 59:33]
  wire  _GEN_208 = _T_67 ? syn[4] : _GEN_138; // @[LTD.scala 55:33]
  wire  syn_new_4 = busy ? syn[4] : _GEN_208; // @[LTD.scala 52:15]
  wire  _GEN_141 = _T_118 ? _GEN_72 : syn[7]; // @[LTD.scala 59:33]
  wire  _GEN_211 = _T_67 ? syn[7] : _GEN_141; // @[LTD.scala 55:33]
  wire  syn_new_7 = busy ? syn[7] : _GEN_211; // @[LTD.scala 52:15]
  wire  _GEN_140 = _T_118 ? _GEN_71 : syn[6]; // @[LTD.scala 59:33]
  wire  _GEN_210 = _T_67 ? syn[6] : _GEN_140; // @[LTD.scala 55:33]
  wire  syn_new_6 = busy ? syn[6] : _GEN_210; // @[LTD.scala 52:15]
  wire [7:0] _T_133 = {syn_new_7,syn_new_6,syn_new_5,syn_new_4,syn_new_3,syn_new_2,syn_new_1,syn_new_0}; // @[LTD.scala 66:40]
  wire  _GEN_143 = _T_118 ? _GEN_74 : syn[9]; // @[LTD.scala 59:33]
  wire  _GEN_213 = _T_67 ? syn[9] : _GEN_143; // @[LTD.scala 55:33]
  wire  syn_new_9 = busy ? syn[9] : _GEN_213; // @[LTD.scala 52:15]
  wire  _GEN_142 = _T_118 ? _GEN_73 : syn[8]; // @[LTD.scala 59:33]
  wire  _GEN_212 = _T_67 ? syn[8] : _GEN_142; // @[LTD.scala 55:33]
  wire  syn_new_8 = busy ? syn[8] : _GEN_212; // @[LTD.scala 52:15]
  wire  _GEN_145 = _T_118 ? _GEN_76 : syn[11]; // @[LTD.scala 59:33]
  wire  _GEN_215 = _T_67 ? syn[11] : _GEN_145; // @[LTD.scala 55:33]
  wire  syn_new_11 = busy ? syn[11] : _GEN_215; // @[LTD.scala 52:15]
  wire  _GEN_144 = _T_118 ? _GEN_75 : syn[10]; // @[LTD.scala 59:33]
  wire  _GEN_214 = _T_67 ? syn[10] : _GEN_144; // @[LTD.scala 55:33]
  wire  syn_new_10 = busy ? syn[10] : _GEN_214; // @[LTD.scala 52:15]
  wire  _GEN_147 = _T_118 ? _GEN_78 : syn[13]; // @[LTD.scala 59:33]
  wire  _GEN_217 = _T_67 ? syn[13] : _GEN_147; // @[LTD.scala 55:33]
  wire  syn_new_13 = busy ? syn[13] : _GEN_217; // @[LTD.scala 52:15]
  wire  _GEN_146 = _T_118 ? _GEN_77 : syn[12]; // @[LTD.scala 59:33]
  wire  _GEN_216 = _T_67 ? syn[12] : _GEN_146; // @[LTD.scala 55:33]
  wire  syn_new_12 = busy ? syn[12] : _GEN_216; // @[LTD.scala 52:15]
  wire  _GEN_149 = _T_118 ? _GEN_80 : syn[15]; // @[LTD.scala 59:33]
  wire  _GEN_219 = _T_67 ? syn[15] : _GEN_149; // @[LTD.scala 55:33]
  wire  syn_new_15 = busy ? syn[15] : _GEN_219; // @[LTD.scala 52:15]
  wire  _GEN_148 = _T_118 ? _GEN_79 : syn[14]; // @[LTD.scala 59:33]
  wire  _GEN_218 = _T_67 ? syn[14] : _GEN_148; // @[LTD.scala 55:33]
  wire  syn_new_14 = busy ? syn[14] : _GEN_218; // @[LTD.scala 52:15]
  wire [15:0] _T_141 = {syn_new_15,syn_new_14,syn_new_13,syn_new_12,syn_new_11,syn_new_10,syn_new_9,syn_new_8,_T_133}; // @[LTD.scala 66:40]
  wire  _GEN_151 = _T_118 ? _GEN_82 : syn[17]; // @[LTD.scala 59:33]
  wire  _GEN_221 = _T_67 ? syn[17] : _GEN_151; // @[LTD.scala 55:33]
  wire  syn_new_17 = busy ? syn[17] : _GEN_221; // @[LTD.scala 52:15]
  wire  _GEN_150 = _T_118 ? _GEN_81 : syn[16]; // @[LTD.scala 59:33]
  wire  _GEN_220 = _T_67 ? syn[16] : _GEN_150; // @[LTD.scala 55:33]
  wire  syn_new_16 = busy ? syn[16] : _GEN_220; // @[LTD.scala 52:15]
  wire  _GEN_153 = _T_118 ? _GEN_84 : syn[19]; // @[LTD.scala 59:33]
  wire  _GEN_223 = _T_67 ? syn[19] : _GEN_153; // @[LTD.scala 55:33]
  wire  syn_new_19 = busy ? syn[19] : _GEN_223; // @[LTD.scala 52:15]
  wire  _GEN_152 = _T_118 ? _GEN_83 : syn[18]; // @[LTD.scala 59:33]
  wire  _GEN_222 = _T_67 ? syn[18] : _GEN_152; // @[LTD.scala 55:33]
  wire  syn_new_18 = busy ? syn[18] : _GEN_222; // @[LTD.scala 52:15]
  wire  _GEN_155 = _T_118 ? _GEN_86 : syn[21]; // @[LTD.scala 59:33]
  wire  _GEN_225 = _T_67 ? syn[21] : _GEN_155; // @[LTD.scala 55:33]
  wire  syn_new_21 = busy ? syn[21] : _GEN_225; // @[LTD.scala 52:15]
  wire  _GEN_154 = _T_118 ? _GEN_85 : syn[20]; // @[LTD.scala 59:33]
  wire  _GEN_224 = _T_67 ? syn[20] : _GEN_154; // @[LTD.scala 55:33]
  wire  syn_new_20 = busy ? syn[20] : _GEN_224; // @[LTD.scala 52:15]
  wire  _GEN_157 = _T_118 ? _GEN_88 : syn[23]; // @[LTD.scala 59:33]
  wire  _GEN_227 = _T_67 ? syn[23] : _GEN_157; // @[LTD.scala 55:33]
  wire  syn_new_23 = busy ? syn[23] : _GEN_227; // @[LTD.scala 52:15]
  wire  _GEN_156 = _T_118 ? _GEN_87 : syn[22]; // @[LTD.scala 59:33]
  wire  _GEN_226 = _T_67 ? syn[22] : _GEN_156; // @[LTD.scala 55:33]
  wire  syn_new_22 = busy ? syn[22] : _GEN_226; // @[LTD.scala 52:15]
  wire [7:0] _T_148 = {syn_new_23,syn_new_22,syn_new_21,syn_new_20,syn_new_19,syn_new_18,syn_new_17,syn_new_16}; // @[LTD.scala 66:40]
  wire  _GEN_159 = _T_118 ? _GEN_90 : syn[25]; // @[LTD.scala 59:33]
  wire  _GEN_229 = _T_67 ? syn[25] : _GEN_159; // @[LTD.scala 55:33]
  wire  syn_new_25 = busy ? syn[25] : _GEN_229; // @[LTD.scala 52:15]
  wire  _GEN_158 = _T_118 ? _GEN_89 : syn[24]; // @[LTD.scala 59:33]
  wire  _GEN_228 = _T_67 ? syn[24] : _GEN_158; // @[LTD.scala 55:33]
  wire  syn_new_24 = busy ? syn[24] : _GEN_228; // @[LTD.scala 52:15]
  wire  _GEN_161 = _T_118 ? _GEN_92 : syn[27]; // @[LTD.scala 59:33]
  wire  _GEN_231 = _T_67 ? syn[27] : _GEN_161; // @[LTD.scala 55:33]
  wire  syn_new_27 = busy ? syn[27] : _GEN_231; // @[LTD.scala 52:15]
  wire  _GEN_160 = _T_118 ? _GEN_91 : syn[26]; // @[LTD.scala 59:33]
  wire  _GEN_230 = _T_67 ? syn[26] : _GEN_160; // @[LTD.scala 55:33]
  wire  syn_new_26 = busy ? syn[26] : _GEN_230; // @[LTD.scala 52:15]
  wire  _GEN_163 = _T_118 ? _GEN_94 : syn[29]; // @[LTD.scala 59:33]
  wire  _GEN_233 = _T_67 ? syn[29] : _GEN_163; // @[LTD.scala 55:33]
  wire  syn_new_29 = busy ? syn[29] : _GEN_233; // @[LTD.scala 52:15]
  wire  _GEN_162 = _T_118 ? _GEN_93 : syn[28]; // @[LTD.scala 59:33]
  wire  _GEN_232 = _T_67 ? syn[28] : _GEN_162; // @[LTD.scala 55:33]
  wire  syn_new_28 = busy ? syn[28] : _GEN_232; // @[LTD.scala 52:15]
  wire  _GEN_165 = _T_118 ? _GEN_96 : syn[31]; // @[LTD.scala 59:33]
  wire  _GEN_235 = _T_67 ? syn[31] : _GEN_165; // @[LTD.scala 55:33]
  wire  syn_new_31 = busy ? syn[31] : _GEN_235; // @[LTD.scala 52:15]
  wire  _GEN_164 = _T_118 ? _GEN_95 : syn[30]; // @[LTD.scala 59:33]
  wire  _GEN_234 = _T_67 ? syn[30] : _GEN_164; // @[LTD.scala 55:33]
  wire  syn_new_30 = busy ? syn[30] : _GEN_234; // @[LTD.scala 52:15]
  wire [31:0] _T_157 = {syn_new_31,syn_new_30,syn_new_29,syn_new_28,syn_new_27,syn_new_26,syn_new_25,syn_new_24,_T_148,_T_141}; // @[LTD.scala 66:40]
  wire  _GEN_167 = _T_118 ? _GEN_98 : syn[33]; // @[LTD.scala 59:33]
  wire  _GEN_237 = _T_67 ? syn[33] : _GEN_167; // @[LTD.scala 55:33]
  wire  syn_new_33 = busy ? syn[33] : _GEN_237; // @[LTD.scala 52:15]
  wire  _GEN_166 = _T_118 ? _GEN_97 : syn[32]; // @[LTD.scala 59:33]
  wire  _GEN_236 = _T_67 ? syn[32] : _GEN_166; // @[LTD.scala 55:33]
  wire  syn_new_32 = busy ? syn[32] : _GEN_236; // @[LTD.scala 52:15]
  wire  _GEN_169 = _T_118 ? _GEN_100 : syn[35]; // @[LTD.scala 59:33]
  wire  _GEN_239 = _T_67 ? syn[35] : _GEN_169; // @[LTD.scala 55:33]
  wire  syn_new_35 = busy ? syn[35] : _GEN_239; // @[LTD.scala 52:15]
  wire  _GEN_168 = _T_118 ? _GEN_99 : syn[34]; // @[LTD.scala 59:33]
  wire  _GEN_238 = _T_67 ? syn[34] : _GEN_168; // @[LTD.scala 55:33]
  wire  syn_new_34 = busy ? syn[34] : _GEN_238; // @[LTD.scala 52:15]
  wire  _GEN_171 = _T_118 ? _GEN_102 : syn[37]; // @[LTD.scala 59:33]
  wire  _GEN_241 = _T_67 ? syn[37] : _GEN_171; // @[LTD.scala 55:33]
  wire  syn_new_37 = busy ? syn[37] : _GEN_241; // @[LTD.scala 52:15]
  wire  _GEN_170 = _T_118 ? _GEN_101 : syn[36]; // @[LTD.scala 59:33]
  wire  _GEN_240 = _T_67 ? syn[36] : _GEN_170; // @[LTD.scala 55:33]
  wire  syn_new_36 = busy ? syn[36] : _GEN_240; // @[LTD.scala 52:15]
  wire  _GEN_173 = _T_118 ? _GEN_104 : syn[39]; // @[LTD.scala 59:33]
  wire  _GEN_243 = _T_67 ? syn[39] : _GEN_173; // @[LTD.scala 55:33]
  wire  syn_new_39 = busy ? syn[39] : _GEN_243; // @[LTD.scala 52:15]
  wire  _GEN_172 = _T_118 ? _GEN_103 : syn[38]; // @[LTD.scala 59:33]
  wire  _GEN_242 = _T_67 ? syn[38] : _GEN_172; // @[LTD.scala 55:33]
  wire  syn_new_38 = busy ? syn[38] : _GEN_242; // @[LTD.scala 52:15]
  wire [7:0] _T_164 = {syn_new_39,syn_new_38,syn_new_37,syn_new_36,syn_new_35,syn_new_34,syn_new_33,syn_new_32}; // @[LTD.scala 66:40]
  wire  _GEN_175 = _T_118 ? _GEN_106 : syn[41]; // @[LTD.scala 59:33]
  wire  _GEN_245 = _T_67 ? syn[41] : _GEN_175; // @[LTD.scala 55:33]
  wire  syn_new_41 = busy ? syn[41] : _GEN_245; // @[LTD.scala 52:15]
  wire  _GEN_174 = _T_118 ? _GEN_105 : syn[40]; // @[LTD.scala 59:33]
  wire  _GEN_244 = _T_67 ? syn[40] : _GEN_174; // @[LTD.scala 55:33]
  wire  syn_new_40 = busy ? syn[40] : _GEN_244; // @[LTD.scala 52:15]
  wire  _GEN_177 = _T_118 ? _GEN_108 : syn[43]; // @[LTD.scala 59:33]
  wire  _GEN_247 = _T_67 ? syn[43] : _GEN_177; // @[LTD.scala 55:33]
  wire  syn_new_43 = busy ? syn[43] : _GEN_247; // @[LTD.scala 52:15]
  wire  _GEN_176 = _T_118 ? _GEN_107 : syn[42]; // @[LTD.scala 59:33]
  wire  _GEN_246 = _T_67 ? syn[42] : _GEN_176; // @[LTD.scala 55:33]
  wire  syn_new_42 = busy ? syn[42] : _GEN_246; // @[LTD.scala 52:15]
  wire  _GEN_179 = _T_118 ? _GEN_110 : syn[45]; // @[LTD.scala 59:33]
  wire  _GEN_249 = _T_67 ? syn[45] : _GEN_179; // @[LTD.scala 55:33]
  wire  syn_new_45 = busy ? syn[45] : _GEN_249; // @[LTD.scala 52:15]
  wire  _GEN_178 = _T_118 ? _GEN_109 : syn[44]; // @[LTD.scala 59:33]
  wire  _GEN_248 = _T_67 ? syn[44] : _GEN_178; // @[LTD.scala 55:33]
  wire  syn_new_44 = busy ? syn[44] : _GEN_248; // @[LTD.scala 52:15]
  wire  _GEN_181 = _T_118 ? _GEN_112 : syn[47]; // @[LTD.scala 59:33]
  wire  _GEN_251 = _T_67 ? syn[47] : _GEN_181; // @[LTD.scala 55:33]
  wire  syn_new_47 = busy ? syn[47] : _GEN_251; // @[LTD.scala 52:15]
  wire  _GEN_180 = _T_118 ? _GEN_111 : syn[46]; // @[LTD.scala 59:33]
  wire  _GEN_250 = _T_67 ? syn[46] : _GEN_180; // @[LTD.scala 55:33]
  wire  syn_new_46 = busy ? syn[46] : _GEN_250; // @[LTD.scala 52:15]
  wire [15:0] _T_172 = {syn_new_47,syn_new_46,syn_new_45,syn_new_44,syn_new_43,syn_new_42,syn_new_41,syn_new_40,_T_164}; // @[LTD.scala 66:40]
  wire  _GEN_183 = _T_118 ? _GEN_114 : syn[49]; // @[LTD.scala 59:33]
  wire  _GEN_253 = _T_67 ? syn[49] : _GEN_183; // @[LTD.scala 55:33]
  wire  syn_new_49 = busy ? syn[49] : _GEN_253; // @[LTD.scala 52:15]
  wire  _GEN_182 = _T_118 ? _GEN_113 : syn[48]; // @[LTD.scala 59:33]
  wire  _GEN_252 = _T_67 ? syn[48] : _GEN_182; // @[LTD.scala 55:33]
  wire  syn_new_48 = busy ? syn[48] : _GEN_252; // @[LTD.scala 52:15]
  wire  _GEN_185 = _T_118 ? _GEN_116 : syn[51]; // @[LTD.scala 59:33]
  wire  _GEN_255 = _T_67 ? syn[51] : _GEN_185; // @[LTD.scala 55:33]
  wire  syn_new_51 = busy ? syn[51] : _GEN_255; // @[LTD.scala 52:15]
  wire  _GEN_184 = _T_118 ? _GEN_115 : syn[50]; // @[LTD.scala 59:33]
  wire  _GEN_254 = _T_67 ? syn[50] : _GEN_184; // @[LTD.scala 55:33]
  wire  syn_new_50 = busy ? syn[50] : _GEN_254; // @[LTD.scala 52:15]
  wire  _GEN_187 = _T_118 ? _GEN_118 : syn[53]; // @[LTD.scala 59:33]
  wire  _GEN_257 = _T_67 ? syn[53] : _GEN_187; // @[LTD.scala 55:33]
  wire  syn_new_53 = busy ? syn[53] : _GEN_257; // @[LTD.scala 52:15]
  wire  _GEN_186 = _T_118 ? _GEN_117 : syn[52]; // @[LTD.scala 59:33]
  wire  _GEN_256 = _T_67 ? syn[52] : _GEN_186; // @[LTD.scala 55:33]
  wire  syn_new_52 = busy ? syn[52] : _GEN_256; // @[LTD.scala 52:15]
  wire  _GEN_189 = _T_118 ? _GEN_120 : syn[55]; // @[LTD.scala 59:33]
  wire  _GEN_259 = _T_67 ? syn[55] : _GEN_189; // @[LTD.scala 55:33]
  wire  syn_new_55 = busy ? syn[55] : _GEN_259; // @[LTD.scala 52:15]
  wire  _GEN_188 = _T_118 ? _GEN_119 : syn[54]; // @[LTD.scala 59:33]
  wire  _GEN_258 = _T_67 ? syn[54] : _GEN_188; // @[LTD.scala 55:33]
  wire  syn_new_54 = busy ? syn[54] : _GEN_258; // @[LTD.scala 52:15]
  wire [7:0] _T_179 = {syn_new_55,syn_new_54,syn_new_53,syn_new_52,syn_new_51,syn_new_50,syn_new_49,syn_new_48}; // @[LTD.scala 66:40]
  wire  _GEN_191 = _T_118 ? _GEN_122 : syn[57]; // @[LTD.scala 59:33]
  wire  _GEN_261 = _T_67 ? syn[57] : _GEN_191; // @[LTD.scala 55:33]
  wire  syn_new_57 = busy ? syn[57] : _GEN_261; // @[LTD.scala 52:15]
  wire  _GEN_190 = _T_118 ? _GEN_121 : syn[56]; // @[LTD.scala 59:33]
  wire  _GEN_260 = _T_67 ? syn[56] : _GEN_190; // @[LTD.scala 55:33]
  wire  syn_new_56 = busy ? syn[56] : _GEN_260; // @[LTD.scala 52:15]
  wire  _GEN_193 = _T_118 ? _GEN_124 : syn[59]; // @[LTD.scala 59:33]
  wire  _GEN_263 = _T_67 ? syn[59] : _GEN_193; // @[LTD.scala 55:33]
  wire  syn_new_59 = busy ? syn[59] : _GEN_263; // @[LTD.scala 52:15]
  wire  _GEN_192 = _T_118 ? _GEN_123 : syn[58]; // @[LTD.scala 59:33]
  wire  _GEN_262 = _T_67 ? syn[58] : _GEN_192; // @[LTD.scala 55:33]
  wire  syn_new_58 = busy ? syn[58] : _GEN_262; // @[LTD.scala 52:15]
  wire  _GEN_195 = _T_118 ? _GEN_126 : syn[61]; // @[LTD.scala 59:33]
  wire  _GEN_265 = _T_67 ? syn[61] : _GEN_195; // @[LTD.scala 55:33]
  wire  syn_new_61 = busy ? syn[61] : _GEN_265; // @[LTD.scala 52:15]
  wire  _GEN_194 = _T_118 ? _GEN_125 : syn[60]; // @[LTD.scala 59:33]
  wire  _GEN_264 = _T_67 ? syn[60] : _GEN_194; // @[LTD.scala 55:33]
  wire  syn_new_60 = busy ? syn[60] : _GEN_264; // @[LTD.scala 52:15]
  wire  _GEN_197 = _T_118 ? _GEN_128 : syn[63]; // @[LTD.scala 59:33]
  wire  _GEN_267 = _T_67 ? syn[63] : _GEN_197; // @[LTD.scala 55:33]
  wire  syn_new_63 = busy ? syn[63] : _GEN_267; // @[LTD.scala 52:15]
  wire  _GEN_196 = _T_118 ? _GEN_127 : syn[62]; // @[LTD.scala 59:33]
  wire  _GEN_266 = _T_67 ? syn[62] : _GEN_196; // @[LTD.scala 55:33]
  wire  syn_new_62 = busy ? syn[62] : _GEN_266; // @[LTD.scala 52:15]
  wire [31:0] _T_188 = {syn_new_63,syn_new_62,syn_new_61,syn_new_60,syn_new_59,syn_new_58,syn_new_57,syn_new_56,_T_179,_T_172}; // @[LTD.scala 66:40]
  wire  _T_191 = state == 2'h3; // @[LTD.scala 68:22]
  MaxPeriodFibonacciLFSR MaxPeriodFibonacciLFSR ( // @[PRNG.scala 82:22]
    .clock(MaxPeriodFibonacciLFSR_clock),
    .reset(MaxPeriodFibonacciLFSR_reset),
    .io_out_0(MaxPeriodFibonacciLFSR_io_out_0),
    .io_out_1(MaxPeriodFibonacciLFSR_io_out_1),
    .io_out_2(MaxPeriodFibonacciLFSR_io_out_2),
    .io_out_3(MaxPeriodFibonacciLFSR_io_out_3),
    .io_out_4(MaxPeriodFibonacciLFSR_io_out_4),
    .io_out_5(MaxPeriodFibonacciLFSR_io_out_5),
    .io_out_6(MaxPeriodFibonacciLFSR_io_out_6),
    .io_out_7(MaxPeriodFibonacciLFSR_io_out_7),
    .io_out_8(MaxPeriodFibonacciLFSR_io_out_8),
    .io_out_9(MaxPeriodFibonacciLFSR_io_out_9),
    .io_out_10(MaxPeriodFibonacciLFSR_io_out_10),
    .io_out_11(MaxPeriodFibonacciLFSR_io_out_11),
    .io_out_12(MaxPeriodFibonacciLFSR_io_out_12),
    .io_out_13(MaxPeriodFibonacciLFSR_io_out_13),
    .io_out_14(MaxPeriodFibonacciLFSR_io_out_14),
    .io_out_15(MaxPeriodFibonacciLFSR_io_out_15)
  );
  assign io_in_ready = state == 2'h0; // @[LTD.scala 73:17]
  assign io_out_valid = state == 2'h3; // @[LTD.scala 74:18]
  assign io_out_bits_res = {_T_188,_T_157}; // @[LTD.scala 70:25]
  assign io_out_bits_ret = {_T_188,_T_157}; // @[LTD.scala 66:29]
  assign io_out_bits_cnt = {{58'd0}, value}; // @[LTD.scala 75:21]
  assign MaxPeriodFibonacciLFSR_clock = clock;
  assign MaxPeriodFibonacciLFSR_reset = reset;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  syn = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  r = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      syn <= 64'h0;
    end else begin
      syn <= io_in_bits_syn;
    end
    if (reset) begin
      r <= 10'h0;
    end else if (!(busy)) begin
      if (_T_67) begin
        r <= _T_117;
      end
    end
    if (reset) begin
      value <= 6'h0;
    end else if (!(busy)) begin
      if (!(_T_67)) begin
        if (_T_118) begin
          value <= _T_125;
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else if (busy) begin
      state <= 2'h1;
    end else if (_T_67) begin
      state <= 2'h2;
    end else if (_T_118) begin
      if (_T_123) begin
        state <= 2'h3;
      end else if (_T_126) begin
        state <= 2'h1;
      end
    end else if (_T_191) begin
      state <= 2'h0;
    end
  end
endmodule
module SNN(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [63:0] io_in_bits_src1,
  input  [63:0] io_in_bits_src2,
  input  [6:0]  io_in_bits_func,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits,
  input  [63:0] io_imm,
  input  [63:0] io_srf_0,
  input  [63:0] io_srf_1,
  input  [63:0] io_srf_2,
  input  [63:0] io_srf_3,
  output [2:0]  io_srfAddrGen,
  output        io_wen
);
  wire  ssp_io_in_valid; // @[SNN.scala 98:21]
  wire [63:0] ssp_io_in_bits_src1; // @[SNN.scala 98:21]
  wire [63:0] ssp_io_in_bits_src2; // @[SNN.scala 98:21]
  wire [63:0] ssp_io_in_bits_op; // @[SNN.scala 98:21]
  wire  ssp_io_out_valid; // @[SNN.scala 98:21]
  wire [63:0] ssp_io_out_bits; // @[SNN.scala 98:21]
  wire  neuron_io_in_valid; // @[SNN.scala 106:24]
  wire [63:0] neuron_io_in_bits_src1; // @[SNN.scala 106:24]
  wire [63:0] neuron_io_in_bits_src2; // @[SNN.scala 106:24]
  wire [63:0] neuron_io_in_bits_vinit; // @[SNN.scala 106:24]
  wire [63:0] neuron_io_in_bits_vleak; // @[SNN.scala 106:24]
  wire [63:0] neuron_io_in_bits_spike; // @[SNN.scala 106:24]
  wire [63:0] neuron_io_in_bits_option; // @[SNN.scala 106:24]
  wire  neuron_io_out_valid; // @[SNN.scala 106:24]
  wire [63:0] neuron_io_out_bits; // @[SNN.scala 106:24]
  wire  stdp_io_in_valid; // @[SNN.scala 119:22]
  wire [63:0] stdp_io_in_bits_src1; // @[SNN.scala 119:22]
  wire [63:0] stdp_io_in_bits_src2; // @[SNN.scala 119:22]
  wire [63:0] stdp_io_in_bits_op; // @[SNN.scala 119:22]
  wire [63:0] stdp_io_in_bits_imm; // @[SNN.scala 119:22]
  wire [63:0] stdp_io_in_bits_output; // @[SNN.scala 119:22]
  wire [63:0] stdp_io_in_bits_vinit; // @[SNN.scala 119:22]
  wire  stdp_io_out_valid; // @[SNN.scala 119:22]
  wire [63:0] stdp_io_out_bits_res; // @[SNN.scala 119:22]
  wire  ltd_clock; // @[SNN.scala 130:21]
  wire  ltd_reset; // @[SNN.scala 130:21]
  wire  ltd_io_in_ready; // @[SNN.scala 130:21]
  wire  ltd_io_in_valid; // @[SNN.scala 130:21]
  wire [63:0] ltd_io_in_bits_prob; // @[SNN.scala 130:21]
  wire [63:0] ltd_io_in_bits_syn; // @[SNN.scala 130:21]
  wire  ltd_io_out_valid; // @[SNN.scala 130:21]
  wire [63:0] ltd_io_out_bits_res; // @[SNN.scala 130:21]
  wire [63:0] ltd_io_out_bits_ret; // @[SNN.scala 130:21]
  wire [63:0] ltd_io_out_bits_cnt; // @[SNN.scala 130:21]
  wire  _T = 7'h0 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_1 = 7'h4 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_2 = 7'h1 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_3 = 7'h9 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_4 = 7'h11 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_5 = 7'h19 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_6 = 7'h2 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_7 = 7'he == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_8 = 7'h21 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_9 = 7'h1e == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire [1:0] _T_14 = _T_4 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_15 = _T_5 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_17 = _T_7 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_18 = _T_8 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_19 = _T_9 ? 2'h3 : 2'h0; // @[Mux.scala 27:72]
  wire  _T_22 = _T_1 | _T_3; // @[Mux.scala 27:72]
  wire [1:0] _GEN_5 = {{1'd0}, _T_22}; // @[Mux.scala 27:72]
  wire [1:0] _T_23 = _GEN_5 | _T_14; // @[Mux.scala 27:72]
  wire [1:0] _T_24 = _T_23 | _T_15; // @[Mux.scala 27:72]
  wire [1:0] _GEN_6 = {{1'd0}, _T_6}; // @[Mux.scala 27:72]
  wire [1:0] _T_25 = _T_24 | _GEN_6; // @[Mux.scala 27:72]
  wire [1:0] _T_26 = _T_25 | _T_17; // @[Mux.scala 27:72]
  wire [1:0] _T_27 = _T_26 | _T_18; // @[Mux.scala 27:72]
  wire [1:0] calcUnit = _T_27 | _T_19; // @[Mux.scala 27:72]
  wire  _T_29 = calcUnit == 2'h0; // @[SNN.scala 103:43]
  wire  _T_31 = calcUnit == 2'h1; // @[SNN.scala 115:51]
  wire  _T_33 = calcUnit == 2'h2; // @[SNN.scala 125:45]
  wire  _T_35 = calcUnit == 2'h3; // @[SNN.scala 132:35]
  wire  _T_37 = ltd_io_out_bits_cnt != 64'h0; // @[SNN.scala 135:35]
  wire [63:0] _T_49 = _T ? ssp_io_out_bits : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_50 = _T_1 ? neuron_io_out_bits : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_51 = _T_2 ? ssp_io_out_bits : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_52 = _T_3 ? neuron_io_out_bits : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_53 = _T_5 ? stdp_io_out_bits_res : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_54 = _T_6 ? neuron_io_out_bits : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_55 = _T_7 ? stdp_io_out_bits_res : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_56 = _T_4 ? stdp_io_out_bits_res : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_57 = _T_8 ? stdp_io_out_bits_res : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_58 = _T_9 ? ltd_io_out_bits_res : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_59 = _T_49 | _T_50; // @[Mux.scala 27:72]
  wire [63:0] _T_60 = _T_59 | _T_51; // @[Mux.scala 27:72]
  wire [63:0] _T_61 = _T_60 | _T_52; // @[Mux.scala 27:72]
  wire [63:0] _T_62 = _T_61 | _T_53; // @[Mux.scala 27:72]
  wire [63:0] _T_63 = _T_62 | _T_54; // @[Mux.scala 27:72]
  wire [63:0] _T_64 = _T_63 | _T_55; // @[Mux.scala 27:72]
  wire [63:0] _T_65 = _T_64 | _T_56; // @[Mux.scala 27:72]
  wire [63:0] _T_66 = _T_65 | _T_57; // @[Mux.scala 27:72]
  wire [1:0] _T_76 = _T_3 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_77 = _T_1 ? 2'h3 : 2'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_78 = _T_5 ? 3'h4 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_79 = _T_9 ? 3'h4 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_81 = _T_8 ? 3'h5 : 3'h0; // @[Mux.scala 27:72]
  wire [1:0] _GEN_7 = {{1'd0}, _T_7}; // @[Mux.scala 27:72]
  wire [1:0] _T_82 = _GEN_7 | _T_76; // @[Mux.scala 27:72]
  wire [1:0] _T_83 = _T_82 | _T_77; // @[Mux.scala 27:72]
  wire [2:0] _GEN_8 = {{1'd0}, _T_83}; // @[Mux.scala 27:72]
  wire [2:0] _T_84 = _GEN_8 | _T_78; // @[Mux.scala 27:72]
  wire [2:0] _T_85 = _T_84 | _T_79; // @[Mux.scala 27:72]
  wire [2:0] _GEN_9 = {{1'd0}, _T_14}; // @[Mux.scala 27:72]
  wire [2:0] _T_86 = _T_85 | _GEN_9; // @[Mux.scala 27:72]
  wire  _T_88 = 2'h0 == calcUnit; // @[LookupTree.scala 24:34]
  wire  _T_89 = 2'h1 == calcUnit; // @[LookupTree.scala 24:34]
  wire  _T_90 = 2'h2 == calcUnit; // @[LookupTree.scala 24:34]
  wire  _T_91 = 2'h3 == calcUnit; // @[LookupTree.scala 24:34]
  wire  _T_100 = io_in_bits_func == 7'h4; // @[SNN.scala 39:41]
  wire  _T_101 = io_in_bits_func == 7'he; // @[SNN.scala 39:57]
  wire  _T_102 = _T_100 | _T_101; // @[SNN.scala 39:49]
  wire  _T_103 = io_in_bits_func == 7'h9; // @[SNN.scala 39:75]
  wire  _T_104 = _T_102 | _T_103; // @[SNN.scala 39:67]
  wire  _T_105 = io_in_bits_func == 7'h19; // @[SNN.scala 39:91]
  wire  _T_106 = _T_104 | _T_105; // @[SNN.scala 39:83]
  wire  _T_107 = io_in_bits_func == 7'h11; // @[SNN.scala 39:107]
  wire  _T_108 = _T_106 | _T_107; // @[SNN.scala 39:99]
  wire  _T_109 = io_in_bits_func == 7'h21; // @[SNN.scala 39:123]
  wire  _T_110 = _T_108 | _T_109; // @[SNN.scala 39:115]
  wire  _T_111 = io_in_bits_func == 7'h1e; // @[SNN.scala 39:141]
  wire  _T_117 = _T_88 & ssp_io_out_valid; // @[Mux.scala 27:72]
  wire  _T_118 = _T_89 & neuron_io_out_valid; // @[Mux.scala 27:72]
  wire  _T_119 = _T_90 & stdp_io_out_valid; // @[Mux.scala 27:72]
  wire  _T_120 = _T_91 & ltd_io_out_valid; // @[Mux.scala 27:72]
  wire  _T_121 = _T_117 | _T_118; // @[Mux.scala 27:72]
  wire  _T_122 = _T_121 | _T_119; // @[Mux.scala 27:72]
  SpikeProc ssp ( // @[SNN.scala 98:21]
    .io_in_valid(ssp_io_in_valid),
    .io_in_bits_src1(ssp_io_in_bits_src1),
    .io_in_bits_src2(ssp_io_in_bits_src2),
    .io_in_bits_op(ssp_io_in_bits_op),
    .io_out_valid(ssp_io_out_valid),
    .io_out_bits(ssp_io_out_bits)
  );
  NeurModule neuron ( // @[SNN.scala 106:24]
    .io_in_valid(neuron_io_in_valid),
    .io_in_bits_src1(neuron_io_in_bits_src1),
    .io_in_bits_src2(neuron_io_in_bits_src2),
    .io_in_bits_vinit(neuron_io_in_bits_vinit),
    .io_in_bits_vleak(neuron_io_in_bits_vleak),
    .io_in_bits_spike(neuron_io_in_bits_spike),
    .io_in_bits_option(neuron_io_in_bits_option),
    .io_out_valid(neuron_io_out_valid),
    .io_out_bits(neuron_io_out_bits)
  );
  STDP stdp ( // @[SNN.scala 119:22]
    .io_in_valid(stdp_io_in_valid),
    .io_in_bits_src1(stdp_io_in_bits_src1),
    .io_in_bits_src2(stdp_io_in_bits_src2),
    .io_in_bits_op(stdp_io_in_bits_op),
    .io_in_bits_imm(stdp_io_in_bits_imm),
    .io_in_bits_output(stdp_io_in_bits_output),
    .io_in_bits_vinit(stdp_io_in_bits_vinit),
    .io_out_valid(stdp_io_out_valid),
    .io_out_bits_res(stdp_io_out_bits_res)
  );
  LTD ltd ( // @[SNN.scala 130:21]
    .clock(ltd_clock),
    .reset(ltd_reset),
    .io_in_ready(ltd_io_in_ready),
    .io_in_valid(ltd_io_in_valid),
    .io_in_bits_prob(ltd_io_in_bits_prob),
    .io_in_bits_syn(ltd_io_in_bits_syn),
    .io_out_valid(ltd_io_out_valid),
    .io_out_bits_res(ltd_io_out_bits_res),
    .io_out_bits_ret(ltd_io_out_bits_ret),
    .io_out_bits_cnt(ltd_io_out_bits_cnt)
  );
  assign io_out_valid = _T_122 | _T_120; // @[SNN.scala 171:18]
  assign io_out_bits = _T_66 | _T_58; // @[SNN.scala 168:17]
  assign io_srfAddrGen = _T_86 | _T_81; // @[SNN.scala 169:19]
  assign io_wen = _T_110 | _T_111; // @[SNN.scala 170:13]
  assign ssp_io_in_valid = io_in_valid & _T_29; // @[SNN.scala 103:21]
  assign ssp_io_in_bits_src1 = io_in_bits_src1; // @[SNN.scala 99:25]
  assign ssp_io_in_bits_src2 = io_in_bits_src2; // @[SNN.scala 100:25]
  assign ssp_io_in_bits_op = {{57'd0}, io_in_bits_func}; // @[SNN.scala 101:23]
  assign neuron_io_in_valid = io_in_valid & _T_31; // @[SNN.scala 115:29]
  assign neuron_io_in_bits_src1 = io_in_bits_src1; // @[SNN.scala 107:29]
  assign neuron_io_in_bits_src2 = io_in_bits_src2; // @[SNN.scala 108:29]
  assign neuron_io_in_bits_vinit = io_srf_1; // @[SNN.scala 110:29]
  assign neuron_io_in_bits_vleak = io_srf_0; // @[SNN.scala 112:29]
  assign neuron_io_in_bits_spike = io_srf_3; // @[SNN.scala 111:29]
  assign neuron_io_in_bits_option = {{57'd0}, io_in_bits_func}; // @[SNN.scala 113:30]
  assign stdp_io_in_valid = io_in_valid & _T_33; // @[SNN.scala 125:22]
  assign stdp_io_in_bits_src1 = io_in_bits_src1; // @[SNN.scala 120:26]
  assign stdp_io_in_bits_src2 = io_in_bits_src2; // @[SNN.scala 121:26]
  assign stdp_io_in_bits_op = {{57'd0}, io_in_bits_func}; // @[SNN.scala 123:24]
  assign stdp_io_in_bits_imm = io_imm; // @[SNN.scala 122:25]
  assign stdp_io_in_bits_output = io_srf_2; // @[SNN.scala 124:28]
  assign stdp_io_in_bits_vinit = io_srf_1; // @[SNN.scala 127:27]
  assign ltd_clock = clock;
  assign ltd_reset = reset;
  assign ltd_io_in_valid = _T_35 & io_in_valid; // @[SNN.scala 132:21]
  assign ltd_io_in_bits_prob = io_in_bits_src1; // @[SNN.scala 131:25]
  assign ltd_io_in_bits_syn = _T_37 ? ltd_io_out_bits_ret : io_in_bits_src2; // @[SNN.scala 135:24]
endmodule
module EXU(
  input         clock,
  input         reset,
  output        io__in_ready,
  input         io__in_valid,
  input  [63:0] io__in_bits_cf_instr,
  input  [38:0] io__in_bits_cf_pc,
  input  [38:0] io__in_bits_cf_pnpc,
  input         io__in_bits_cf_exceptionVec_1,
  input         io__in_bits_cf_exceptionVec_2,
  input         io__in_bits_cf_exceptionVec_12,
  input         io__in_bits_cf_intrVec_0,
  input         io__in_bits_cf_intrVec_1,
  input         io__in_bits_cf_intrVec_2,
  input         io__in_bits_cf_intrVec_3,
  input         io__in_bits_cf_intrVec_4,
  input         io__in_bits_cf_intrVec_5,
  input         io__in_bits_cf_intrVec_6,
  input         io__in_bits_cf_intrVec_7,
  input         io__in_bits_cf_intrVec_8,
  input         io__in_bits_cf_intrVec_9,
  input         io__in_bits_cf_intrVec_10,
  input         io__in_bits_cf_intrVec_11,
  input  [3:0]  io__in_bits_cf_brIdx,
  input         io__in_bits_cf_crossPageIPFFix,
  input  [2:0]  io__in_bits_ctrl_fuType,
  input  [6:0]  io__in_bits_ctrl_fuOpType,
  input         io__in_bits_ctrl_rfWen,
  input  [4:0]  io__in_bits_ctrl_rfDest,
  input         io__in_bits_ctrl_isNutCoreTrap,
  input  [63:0] io__in_bits_data_src1,
  input  [63:0] io__in_bits_data_src2,
  input  [63:0] io__in_bits_data_imm,
  input  [63:0] io__in_bits_data_srf_0,
  input  [63:0] io__in_bits_data_srf_1,
  input  [63:0] io__in_bits_data_srf_2,
  input  [63:0] io__in_bits_data_srf_3,
  input         io__out_ready,
  output        io__out_valid,
  output [63:0] io__out_bits_decode_cf_instr,
  output [38:0] io__out_bits_decode_cf_pc,
  output [38:0] io__out_bits_decode_cf_redirect_target,
  output        io__out_bits_decode_cf_redirect_valid,
  output [2:0]  io__out_bits_decode_ctrl_fuType,
  output        io__out_bits_decode_ctrl_rfWen,
  output [4:0]  io__out_bits_decode_ctrl_rfDest,
  output        io__out_bits_decode_ctrl_srfWen,
  output [2:0]  io__out_bits_decode_ctrl_srfDest,
  output        io__out_bits_isMMIO,
  output [63:0] io__out_bits_intrNO,
  output [63:0] io__out_bits_commits_0,
  output [63:0] io__out_bits_commits_1,
  output [63:0] io__out_bits_commits_2,
  output [63:0] io__out_bits_commits_3,
  output [63:0] io__out_bits_commits_5,
  input         io__flush,
  input         io__dmem_req_ready,
  output        io__dmem_req_valid,
  output [38:0] io__dmem_req_bits_addr,
  output [2:0]  io__dmem_req_bits_size,
  output [3:0]  io__dmem_req_bits_cmd,
  output [7:0]  io__dmem_req_bits_wmask,
  output [63:0] io__dmem_req_bits_wdata,
  input         io__dmem_resp_valid,
  input  [63:0] io__dmem_resp_bits_rdata,
  output        io__forward_valid,
  output        io__forward_wb_rfWen,
  output [4:0]  io__forward_wb_rfDest,
  output [63:0] io__forward_wb_rfData,
  output [2:0]  io__forward_wb_srfDest,
  output [63:0] io__forward_wb_srfData,
  output [2:0]  io__forward_fuType,
  output [1:0]  io__memMMU_imem_priviledgeMode,
  output [1:0]  io__memMMU_dmem_priviledgeMode,
  output        io__memMMU_dmem_status_sum,
  output        io__memMMU_dmem_status_mxr,
  input         io__memMMU_dmem_loadPF,
  input         io__memMMU_dmem_storePF,
  input  [38:0] io__memMMU_dmem_addr,
  output [63:0] _T_4181,
  output [63:0] _T_4184,
  input         _T_183,
  input         _T_38_0,
  output        flushICache,
  output [63:0] _T_4185,
  output [63:0] satp,
  output        _T_243_valid,
  output [38:0] _T_243_pc,
  output        _T_243_isMissPredict,
  output [38:0] _T_243_actualTarget,
  output        _T_243_actualTaken,
  output [6:0]  _T_243_fuOpType,
  output [1:0]  _T_243_btbType,
  output        _T_243_isRVC,
  output [1:0]  _T_4178,
  input         io_in_valid,
  input         mmio,
  input         _T_186,
  input         io_extra_mtip,
  output        amoReq,
  input         DISPLAY_ENABLE,
  input         io_extra_meip_0,
  input         _T_187,
  input         vmEnable,
  output [11:0] intrVec,
  input         _T_37_1,
  input         io_extra_msip,
  input         _T_65_0,
  output [63:0] _T_4183,
  output [63:0] _T_4182,
  output        flushTLB,
  input         _T_66_0,
  output [63:0] _T_4179,
  input         falseWire_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  alu_clock; // @[EXU.scala 45:19]
  wire  alu_reset; // @[EXU.scala 45:19]
  wire  alu_io_in_valid; // @[EXU.scala 45:19]
  wire [63:0] alu_io_in_bits_src1; // @[EXU.scala 45:19]
  wire [63:0] alu_io_in_bits_src2; // @[EXU.scala 45:19]
  wire [6:0] alu_io_in_bits_func; // @[EXU.scala 45:19]
  wire  alu_io_out_ready; // @[EXU.scala 45:19]
  wire  alu_io_out_valid; // @[EXU.scala 45:19]
  wire [63:0] alu_io_out_bits; // @[EXU.scala 45:19]
  wire [63:0] alu_io_cfIn_instr; // @[EXU.scala 45:19]
  wire [38:0] alu_io_cfIn_pc; // @[EXU.scala 45:19]
  wire [38:0] alu_io_cfIn_pnpc; // @[EXU.scala 45:19]
  wire [3:0] alu_io_cfIn_brIdx; // @[EXU.scala 45:19]
  wire [38:0] alu_io_redirect_target; // @[EXU.scala 45:19]
  wire  alu_io_redirect_valid; // @[EXU.scala 45:19]
  wire [63:0] alu_io_offset; // @[EXU.scala 45:19]
  wire  alu__T_272_0; // @[EXU.scala 45:19]
  wire  alu__T_288_0; // @[EXU.scala 45:19]
  wire  alu__T_308_0; // @[EXU.scala 45:19]
  wire  alu__T_243_0_valid; // @[EXU.scala 45:19]
  wire [38:0] alu__T_243_0_pc; // @[EXU.scala 45:19]
  wire  alu__T_243_0_isMissPredict; // @[EXU.scala 45:19]
  wire [38:0] alu__T_243_0_actualTarget; // @[EXU.scala 45:19]
  wire  alu__T_243_0_actualTaken; // @[EXU.scala 45:19]
  wire [6:0] alu__T_243_0_fuOpType; // @[EXU.scala 45:19]
  wire [1:0] alu__T_243_0_btbType; // @[EXU.scala 45:19]
  wire  alu__T_243_0_isRVC; // @[EXU.scala 45:19]
  wire  alu__T_283_0; // @[EXU.scala 45:19]
  wire  alu__T_249_0; // @[EXU.scala 45:19]
  wire  alu__T_266_0; // @[EXU.scala 45:19]
  wire  alu_DISPLAY_ENABLE; // @[EXU.scala 45:19]
  wire  alu__T_250_1; // @[EXU.scala 45:19]
  wire  alu__T_310_0; // @[EXU.scala 45:19]
  wire  alu__T_304_0; // @[EXU.scala 45:19]
  wire  alu__T_277_0; // @[EXU.scala 45:19]
  wire  alu__T_298_0; // @[EXU.scala 45:19]
  wire  alu__T_294_0; // @[EXU.scala 45:19]
  wire  alu__T_261_0; // @[EXU.scala 45:19]
  wire  alu__T_306_0; // @[EXU.scala 45:19]
  wire  alu__T_255_0; // @[EXU.scala 45:19]
  wire  alu__T_302_0; // @[EXU.scala 45:19]
  wire  lsu_clock; // @[EXU.scala 53:19]
  wire  lsu_reset; // @[EXU.scala 53:19]
  wire  lsu_io__in_ready; // @[EXU.scala 53:19]
  wire  lsu_io__in_valid; // @[EXU.scala 53:19]
  wire [63:0] lsu_io__in_bits_src1; // @[EXU.scala 53:19]
  wire [63:0] lsu_io__in_bits_src2; // @[EXU.scala 53:19]
  wire [6:0] lsu_io__in_bits_func; // @[EXU.scala 53:19]
  wire  lsu_io__out_ready; // @[EXU.scala 53:19]
  wire  lsu_io__out_valid; // @[EXU.scala 53:19]
  wire [63:0] lsu_io__out_bits; // @[EXU.scala 53:19]
  wire [63:0] lsu_io__wdata; // @[EXU.scala 53:19]
  wire [31:0] lsu_io__instr; // @[EXU.scala 53:19]
  wire  lsu_io__dmem_req_ready; // @[EXU.scala 53:19]
  wire  lsu_io__dmem_req_valid; // @[EXU.scala 53:19]
  wire [38:0] lsu_io__dmem_req_bits_addr; // @[EXU.scala 53:19]
  wire [2:0] lsu_io__dmem_req_bits_size; // @[EXU.scala 53:19]
  wire [3:0] lsu_io__dmem_req_bits_cmd; // @[EXU.scala 53:19]
  wire [7:0] lsu_io__dmem_req_bits_wmask; // @[EXU.scala 53:19]
  wire [63:0] lsu_io__dmem_req_bits_wdata; // @[EXU.scala 53:19]
  wire  lsu_io__dmem_resp_valid; // @[EXU.scala 53:19]
  wire [63:0] lsu_io__dmem_resp_bits_rdata; // @[EXU.scala 53:19]
  wire  lsu_io__isMMIO; // @[EXU.scala 53:19]
  wire  lsu_io__dtlbPF; // @[EXU.scala 53:19]
  wire  lsu_io__loadAddrMisaligned; // @[EXU.scala 53:19]
  wire  lsu_io__storeAddrMisaligned; // @[EXU.scala 53:19]
  wire  lsu__T_250; // @[EXU.scala 53:19]
  wire  lsu_setLr_0; // @[EXU.scala 53:19]
  wire  lsu_DTLBPF; // @[EXU.scala 53:19]
  wire  lsu_lsuMMIO_0; // @[EXU.scala 53:19]
  wire  lsu_amoReq_0; // @[EXU.scala 53:19]
  wire  lsu_DISPLAY_ENABLE; // @[EXU.scala 53:19]
  wire  lsu_DTLBENABLE; // @[EXU.scala 53:19]
  wire [63:0] lsu_io_in_bits_src1; // @[EXU.scala 53:19]
  wire  lsu_DTLBFINISH; // @[EXU.scala 53:19]
  wire  lsu__T_258; // @[EXU.scala 53:19]
  wire [63:0] lsu_setLrAddr_0; // @[EXU.scala 53:19]
  wire  lsu__T_262; // @[EXU.scala 53:19]
  wire  lsu_io_isMMIO; // @[EXU.scala 53:19]
  wire  lsu_setLrVal_0; // @[EXU.scala 53:19]
  wire [63:0] lsu_lr_addr; // @[EXU.scala 53:19]
  wire  mdu_clock; // @[EXU.scala 62:19]
  wire  mdu_reset; // @[EXU.scala 62:19]
  wire  mdu_io_in_ready; // @[EXU.scala 62:19]
  wire  mdu_io_in_valid; // @[EXU.scala 62:19]
  wire [63:0] mdu_io_in_bits_src1; // @[EXU.scala 62:19]
  wire [63:0] mdu_io_in_bits_src2; // @[EXU.scala 62:19]
  wire [6:0] mdu_io_in_bits_func; // @[EXU.scala 62:19]
  wire  mdu_io_out_ready; // @[EXU.scala 62:19]
  wire  mdu_io_out_valid; // @[EXU.scala 62:19]
  wire [63:0] mdu_io_out_bits; // @[EXU.scala 62:19]
  wire  mdu_DISPLAY_ENABLE; // @[EXU.scala 62:19]
  wire  mdu__T_87_0; // @[EXU.scala 62:19]
  wire  csr_clock; // @[EXU.scala 67:19]
  wire  csr_reset; // @[EXU.scala 67:19]
  wire  csr_io_in_valid; // @[EXU.scala 67:19]
  wire [63:0] csr_io_in_bits_src1; // @[EXU.scala 67:19]
  wire [63:0] csr_io_in_bits_src2; // @[EXU.scala 67:19]
  wire [6:0] csr_io_in_bits_func; // @[EXU.scala 67:19]
  wire  csr_io_out_ready; // @[EXU.scala 67:19]
  wire  csr_io_out_valid; // @[EXU.scala 67:19]
  wire [63:0] csr_io_out_bits; // @[EXU.scala 67:19]
  wire [63:0] csr_io_cfIn_instr; // @[EXU.scala 67:19]
  wire [38:0] csr_io_cfIn_pc; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_exceptionVec_1; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_exceptionVec_2; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_exceptionVec_4; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_exceptionVec_6; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_exceptionVec_12; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_intrVec_0; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_intrVec_1; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_intrVec_2; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_intrVec_3; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_intrVec_4; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_intrVec_5; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_intrVec_6; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_intrVec_7; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_intrVec_8; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_intrVec_9; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_intrVec_10; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_intrVec_11; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_crossPageIPFFix; // @[EXU.scala 67:19]
  wire [38:0] csr_io_redirect_target; // @[EXU.scala 67:19]
  wire  csr_io_redirect_valid; // @[EXU.scala 67:19]
  wire  csr_io_instrValid; // @[EXU.scala 67:19]
  wire [63:0] csr_io_intrNO; // @[EXU.scala 67:19]
  wire [1:0] csr_io_imemMMU_priviledgeMode; // @[EXU.scala 67:19]
  wire [1:0] csr_io_dmemMMU_priviledgeMode; // @[EXU.scala 67:19]
  wire  csr_io_dmemMMU_status_sum; // @[EXU.scala 67:19]
  wire  csr_io_dmemMMU_status_mxr; // @[EXU.scala 67:19]
  wire  csr_io_dmemMMU_loadPF; // @[EXU.scala 67:19]
  wire  csr_io_dmemMMU_storePF; // @[EXU.scala 67:19]
  wire [38:0] csr_io_dmemMMU_addr; // @[EXU.scala 67:19]
  wire  csr_io_wenFix; // @[EXU.scala 67:19]
  wire [63:0] csr__T_4181_0; // @[EXU.scala 67:19]
  wire  csr_perfCntCondMloadInstr; // @[EXU.scala 67:19]
  wire [63:0] csr__T_4184_0; // @[EXU.scala 67:19]
  wire  csr_perfCntCondMlsuInstr; // @[EXU.scala 67:19]
  wire  csr_set_lr; // @[EXU.scala 67:19]
  wire  csr_perfCntCondMrawStall; // @[EXU.scala 67:19]
  wire  csr_Custom4; // @[EXU.scala 67:19]
  wire  csr_Custom7; // @[EXU.scala 67:19]
  wire [63:0] csr__T_4185_0; // @[EXU.scala 67:19]
  wire  csr_MbpRRight; // @[EXU.scala 67:19]
  wire [63:0] csr_perfCnts_2_0; // @[EXU.scala 67:19]
  wire [63:0] csr_satp_0; // @[EXU.scala 67:19]
  wire [1:0] csr__T_4178_0; // @[EXU.scala 67:19]
  wire  csr_Custom6; // @[EXU.scala 67:19]
  wire  csr_perfCntCondMinstret; // @[EXU.scala 67:19]
  wire  csr_MbpBRight; // @[EXU.scala 67:19]
  wire  csr_perfCntCondMexuBusy; // @[EXU.scala 67:19]
  wire  csr_perfCntCondMmduInstr; // @[EXU.scala 67:19]
  wire  csr_mtip_0; // @[EXU.scala 67:19]
  wire  csr_Custom3; // @[EXU.scala 67:19]
  wire  csr_DISPLAY_ENABLE; // @[EXU.scala 67:19]
  wire  csr_MbpBWrong; // @[EXU.scala 67:19]
  wire  csr_MbpRWrong; // @[EXU.scala 67:19]
  wire  csr_meip_0; // @[EXU.scala 67:19]
  wire  csr_perfCntCondISUIssue; // @[EXU.scala 67:19]
  wire  csr_nutcoretrap_0; // @[EXU.scala 67:19]
  wire  csr_MbpIRight; // @[EXU.scala 67:19]
  wire  csr_perfCntCondMcsrInstr; // @[EXU.scala 67:19]
  wire  csr_perfCntCondMsnnInstr; // @[EXU.scala 67:19]
  wire  csr_perfCntCondMmulInstr; // @[EXU.scala 67:19]
  wire [63:0] csr_LSUADDR; // @[EXU.scala 67:19]
  wire  csr_Custom5; // @[EXU.scala 67:19]
  wire  csr_MbpJRight; // @[EXU.scala 67:19]
  wire  csr_perfCntCondMbruInstr; // @[EXU.scala 67:19]
  wire [11:0] csr_intrVec_0; // @[EXU.scala 67:19]
  wire  csr_perfCntCondMaluInstr; // @[EXU.scala 67:19]
  wire  csr_Custom8; // @[EXU.scala 67:19]
  wire  csr_perfCntCondMloadStall; // @[EXU.scala 67:19]
  wire  csr_Custom2; // @[EXU.scala 67:19]
  wire  csr_msip_0; // @[EXU.scala 67:19]
  wire  csr_MbpIWrong; // @[EXU.scala 67:19]
  wire [63:0] csr_set_lr_addr; // @[EXU.scala 67:19]
  wire  csr_perfCntCondMimemStall; // @[EXU.scala 67:19]
  wire  csr_perfCntCondMstoreStall; // @[EXU.scala 67:19]
  wire [63:0] csr__T_4183_0; // @[EXU.scala 67:19]
  wire [63:0] csr__T_4182_0; // @[EXU.scala 67:19]
  wire [63:0] csr_perfCnts_0_0; // @[EXU.scala 67:19]
  wire  csr_perfCntCondMifuFlush; // @[EXU.scala 67:19]
  wire [63:0] csr__T_4179_0; // @[EXU.scala 67:19]
  wire  csr_perfCntCondMmmioInstr; // @[EXU.scala 67:19]
  wire  csr_perfCntCondMultiCommit; // @[EXU.scala 67:19]
  wire  csr_Custom1; // @[EXU.scala 67:19]
  wire  csr_MbpJWrong; // @[EXU.scala 67:19]
  wire  csr_set_lr_val; // @[EXU.scala 67:19]
  wire [63:0] csr_lrAddr_0; // @[EXU.scala 67:19]
  wire  mou_clock; // @[EXU.scala 81:19]
  wire  mou_reset; // @[EXU.scala 81:19]
  wire  mou_io_in_valid; // @[EXU.scala 81:19]
  wire [6:0] mou_io_in_bits_func; // @[EXU.scala 81:19]
  wire [38:0] mou_io_cfIn_pc; // @[EXU.scala 81:19]
  wire [38:0] mou_io_redirect_target; // @[EXU.scala 81:19]
  wire  mou_io_redirect_valid; // @[EXU.scala 81:19]
  wire  mou_flushICache_0; // @[EXU.scala 81:19]
  wire  mou_DISPLAY_ENABLE; // @[EXU.scala 81:19]
  wire  mou_flushTLB_0; // @[EXU.scala 81:19]
  wire  snn_clock; // @[EXU.scala 87:19]
  wire  snn_reset; // @[EXU.scala 87:19]
  wire  snn_io_in_valid; // @[EXU.scala 87:19]
  wire [63:0] snn_io_in_bits_src1; // @[EXU.scala 87:19]
  wire [63:0] snn_io_in_bits_src2; // @[EXU.scala 87:19]
  wire [6:0] snn_io_in_bits_func; // @[EXU.scala 87:19]
  wire  snn_io_out_ready; // @[EXU.scala 87:19]
  wire  snn_io_out_valid; // @[EXU.scala 87:19]
  wire [63:0] snn_io_out_bits; // @[EXU.scala 87:19]
  wire [63:0] snn_io_imm; // @[EXU.scala 87:19]
  wire [63:0] snn_io_srf_0; // @[EXU.scala 87:19]
  wire [63:0] snn_io_srf_1; // @[EXU.scala 87:19]
  wire [63:0] snn_io_srf_2; // @[EXU.scala 87:19]
  wire [63:0] snn_io_srf_3; // @[EXU.scala 87:19]
  wire [2:0] snn_io_srfAddrGen; // @[EXU.scala 87:19]
  wire  snn_io_wen; // @[EXU.scala 87:19]
  wire  Monitor_clk; // @[EXU.scala 144:21]
  wire  Monitor_reset; // @[EXU.scala 144:21]
  wire  Monitor_isNutCoreTrap; // @[EXU.scala 144:21]
  wire [31:0] Monitor_trapCode; // @[EXU.scala 144:21]
  wire [63:0] Monitor_trapPC; // @[EXU.scala 144:21]
  wire [63:0] Monitor_cycleCnt; // @[EXU.scala 144:21]
  wire [63:0] Monitor_instrCnt; // @[EXU.scala 144:21]
  wire  _T = io__in_bits_ctrl_fuType == 3'h0; // @[EXU.scala 43:57]
  wire  _T_1 = _T & io__in_valid; // @[EXU.scala 43:66]
  wire  _T_2 = ~io__flush; // @[EXU.scala 43:84]
  wire  fuValids_0 = _T_1 & _T_2; // @[EXU.scala 43:81]
  wire  _T_4 = io__in_bits_ctrl_fuType == 3'h1; // @[EXU.scala 43:57]
  wire  _T_5 = _T_4 & io__in_valid; // @[EXU.scala 43:66]
  wire  fuValids_1 = _T_5 & _T_2; // @[EXU.scala 43:81]
  wire  _T_8 = io__in_bits_ctrl_fuType == 3'h2; // @[EXU.scala 43:57]
  wire  _T_9 = _T_8 & io__in_valid; // @[EXU.scala 43:66]
  wire  _T_12 = io__in_bits_ctrl_fuType == 3'h3; // @[EXU.scala 43:57]
  wire  _T_13 = _T_12 & io__in_valid; // @[EXU.scala 43:66]
  wire  fuValids_3 = _T_13 & _T_2; // @[EXU.scala 43:81]
  wire  _T_16 = io__in_bits_ctrl_fuType == 3'h4; // @[EXU.scala 43:57]
  wire  _T_17 = _T_16 & io__in_valid; // @[EXU.scala 43:66]
  wire  _T_20 = io__in_bits_ctrl_fuType == 3'h5; // @[EXU.scala 43:57]
  wire  _T_21 = _T_20 & io__in_valid; // @[EXU.scala 43:66]
  wire [38:0] _T_24 = io__in_bits_cf_pc ^ 39'h30000000; // @[NutCore.scala 86:11]
  wire  _T_26 = _T_24[31:28] == 4'h0; // @[NutCore.scala 86:44]
  wire [38:0] _T_27 = io__in_bits_cf_pc ^ 39'h40000000; // @[NutCore.scala 86:11]
  wire  _T_29 = _T_27[31:30] == 2'h0; // @[NutCore.scala 86:44]
  wire  _T_30 = _T_26 | _T_29; // @[NutCore.scala 87:15]
  wire  _T_31 = _T_30 & io__out_valid; // @[EXU.scala 58:81]
  wire  lsuTlbPF = lsu_io__dtlbPF; // @[UnpipelinedLSU.scala 44:12]
  wire  _T_35 = ~lsuTlbPF; // @[EXU.scala 95:28]
  wire  _T_36 = ~lsu_io__loadAddrMisaligned; // @[EXU.scala 95:41]
  wire  _T_37 = _T_35 & _T_36; // @[EXU.scala 95:38]
  wire  _T_38 = ~lsu_io__storeAddrMisaligned; // @[EXU.scala 95:71]
  wire  _T_39 = _T_37 & _T_38; // @[EXU.scala 95:68]
  wire  _T_40 = ~fuValids_1; // @[EXU.scala 95:102]
  wire  _T_41 = _T_39 | _T_40; // @[EXU.scala 95:99]
  wire  _T_42 = io__in_bits_ctrl_rfWen & _T_41; // @[EXU.scala 95:24]
  wire  _T_43 = csr_io_wenFix & fuValids_3; // @[EXU.scala 95:144]
  wire  _T_44 = ~_T_43; // @[EXU.scala 95:128]
  wire  _T_46 = ~fuValids_0; // @[EXU.scala 98:32]
  wire [38:0] _T_48_target = csr_io_redirect_valid ? csr_io_redirect_target : alu_io_redirect_target; // @[EXU.scala 105:10]
  wire  _T_48_valid = csr_io_redirect_valid ? csr_io_redirect_valid : alu_io_redirect_valid; // @[EXU.scala 105:10]
  wire  _T_50 = mou_io_redirect_valid | csr_io_redirect_valid; // @[EXU.scala 107:31]
  wire  _T_51 = _T_50 | alu_io_redirect_valid; // @[EXU.scala 107:56]
  reg [63:0] _T_52; // @[GTimer.scala 24:20]
  wire [63:0] _T_54 = _T_52 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_56 = _T_51 & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  wire  _T_58 = ~reset; // @[Debug.scala 56:24]
  reg [63:0] _T_63; // @[GTimer.scala 24:20]
  wire [63:0] _T_65 = _T_63 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_72 = 3'h1 == io__in_bits_ctrl_fuType; // @[Mux.scala 80:60]
  wire  _T_73 = _T_72 ? lsu_io__out_valid : 1'h1; // @[Mux.scala 80:57]
  wire  _T_74 = 3'h2 == io__in_bits_ctrl_fuType; // @[Mux.scala 80:60]
  wire  _T_75 = _T_74 ? mdu_io_out_valid : _T_73; // @[Mux.scala 80:57]
  wire  _T_76 = 3'h5 == io__in_bits_ctrl_fuType; // @[Mux.scala 80:60]
  wire  _T_77 = _T_76 ? snn_io_out_valid : _T_75; // @[Mux.scala 80:57]
  wire  _T_79 = ~io__in_valid; // @[EXU.scala 124:18]
  wire  _T_82 = alu_io_out_ready & alu_io_out_valid; // @[Decoupled.scala 40:37]
  wire  isBru = io__in_bits_ctrl_fuOpType[4]; // @[ALU.scala 61:31]
  wire  _T_85 = ~isBru; // @[EXU.scala 136:46]
  wire  _T_86 = _T_82 & _T_85; // @[EXU.scala 136:43]
  wire  _T_88 = _T_82 & isBru; // @[EXU.scala 137:43]
  wire  _T_89 = lsu_io__out_ready & lsu_io__out_valid; // @[Decoupled.scala 40:37]
  wire  _T_90 = mdu_io_out_ready & mdu_io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_91 = snn_io_out_ready & snn_io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_92 = csr_io_out_ready & csr_io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_95 = io__in_bits_ctrl_isNutCoreTrap & io__in_valid; // @[EXU.scala 147:53]
  ALU alu ( // @[EXU.scala 45:19]
    .clock(alu_clock),
    .reset(alu_reset),
    .io_in_valid(alu_io_in_valid),
    .io_in_bits_src1(alu_io_in_bits_src1),
    .io_in_bits_src2(alu_io_in_bits_src2),
    .io_in_bits_func(alu_io_in_bits_func),
    .io_out_ready(alu_io_out_ready),
    .io_out_valid(alu_io_out_valid),
    .io_out_bits(alu_io_out_bits),
    .io_cfIn_instr(alu_io_cfIn_instr),
    .io_cfIn_pc(alu_io_cfIn_pc),
    .io_cfIn_pnpc(alu_io_cfIn_pnpc),
    .io_cfIn_brIdx(alu_io_cfIn_brIdx),
    .io_redirect_target(alu_io_redirect_target),
    .io_redirect_valid(alu_io_redirect_valid),
    .io_offset(alu_io_offset),
    ._T_272_0(alu__T_272_0),
    ._T_288_0(alu__T_288_0),
    ._T_308_0(alu__T_308_0),
    ._T_243_0_valid(alu__T_243_0_valid),
    ._T_243_0_pc(alu__T_243_0_pc),
    ._T_243_0_isMissPredict(alu__T_243_0_isMissPredict),
    ._T_243_0_actualTarget(alu__T_243_0_actualTarget),
    ._T_243_0_actualTaken(alu__T_243_0_actualTaken),
    ._T_243_0_fuOpType(alu__T_243_0_fuOpType),
    ._T_243_0_btbType(alu__T_243_0_btbType),
    ._T_243_0_isRVC(alu__T_243_0_isRVC),
    ._T_283_0(alu__T_283_0),
    ._T_249_0(alu__T_249_0),
    ._T_266_0(alu__T_266_0),
    .DISPLAY_ENABLE(alu_DISPLAY_ENABLE),
    ._T_250_1(alu__T_250_1),
    ._T_310_0(alu__T_310_0),
    ._T_304_0(alu__T_304_0),
    ._T_277_0(alu__T_277_0),
    ._T_298_0(alu__T_298_0),
    ._T_294_0(alu__T_294_0),
    ._T_261_0(alu__T_261_0),
    ._T_306_0(alu__T_306_0),
    ._T_255_0(alu__T_255_0),
    ._T_302_0(alu__T_302_0)
  );
  UnpipelinedLSU lsu ( // @[EXU.scala 53:19]
    .clock(lsu_clock),
    .reset(lsu_reset),
    .io__in_ready(lsu_io__in_ready),
    .io__in_valid(lsu_io__in_valid),
    .io__in_bits_src1(lsu_io__in_bits_src1),
    .io__in_bits_src2(lsu_io__in_bits_src2),
    .io__in_bits_func(lsu_io__in_bits_func),
    .io__out_ready(lsu_io__out_ready),
    .io__out_valid(lsu_io__out_valid),
    .io__out_bits(lsu_io__out_bits),
    .io__wdata(lsu_io__wdata),
    .io__instr(lsu_io__instr),
    .io__dmem_req_ready(lsu_io__dmem_req_ready),
    .io__dmem_req_valid(lsu_io__dmem_req_valid),
    .io__dmem_req_bits_addr(lsu_io__dmem_req_bits_addr),
    .io__dmem_req_bits_size(lsu_io__dmem_req_bits_size),
    .io__dmem_req_bits_cmd(lsu_io__dmem_req_bits_cmd),
    .io__dmem_req_bits_wmask(lsu_io__dmem_req_bits_wmask),
    .io__dmem_req_bits_wdata(lsu_io__dmem_req_bits_wdata),
    .io__dmem_resp_valid(lsu_io__dmem_resp_valid),
    .io__dmem_resp_bits_rdata(lsu_io__dmem_resp_bits_rdata),
    .io__isMMIO(lsu_io__isMMIO),
    .io__dtlbPF(lsu_io__dtlbPF),
    .io__loadAddrMisaligned(lsu_io__loadAddrMisaligned),
    .io__storeAddrMisaligned(lsu_io__storeAddrMisaligned),
    ._T_250(lsu__T_250),
    .setLr_0(lsu_setLr_0),
    .DTLBPF(lsu_DTLBPF),
    .lsuMMIO_0(lsu_lsuMMIO_0),
    .amoReq_0(lsu_amoReq_0),
    .DISPLAY_ENABLE(lsu_DISPLAY_ENABLE),
    .DTLBENABLE(lsu_DTLBENABLE),
    .io_in_bits_src1(lsu_io_in_bits_src1),
    .DTLBFINISH(lsu_DTLBFINISH),
    ._T_258(lsu__T_258),
    .setLrAddr_0(lsu_setLrAddr_0),
    ._T_262(lsu__T_262),
    .io_isMMIO(lsu_io_isMMIO),
    .setLrVal_0(lsu_setLrVal_0),
    .lr_addr(lsu_lr_addr)
  );
  MDU mdu ( // @[EXU.scala 62:19]
    .clock(mdu_clock),
    .reset(mdu_reset),
    .io_in_ready(mdu_io_in_ready),
    .io_in_valid(mdu_io_in_valid),
    .io_in_bits_src1(mdu_io_in_bits_src1),
    .io_in_bits_src2(mdu_io_in_bits_src2),
    .io_in_bits_func(mdu_io_in_bits_func),
    .io_out_ready(mdu_io_out_ready),
    .io_out_valid(mdu_io_out_valid),
    .io_out_bits(mdu_io_out_bits),
    .DISPLAY_ENABLE(mdu_DISPLAY_ENABLE),
    ._T_87_0(mdu__T_87_0)
  );
  CSR csr ( // @[EXU.scala 67:19]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_in_valid(csr_io_in_valid),
    .io_in_bits_src1(csr_io_in_bits_src1),
    .io_in_bits_src2(csr_io_in_bits_src2),
    .io_in_bits_func(csr_io_in_bits_func),
    .io_out_ready(csr_io_out_ready),
    .io_out_valid(csr_io_out_valid),
    .io_out_bits(csr_io_out_bits),
    .io_cfIn_instr(csr_io_cfIn_instr),
    .io_cfIn_pc(csr_io_cfIn_pc),
    .io_cfIn_exceptionVec_1(csr_io_cfIn_exceptionVec_1),
    .io_cfIn_exceptionVec_2(csr_io_cfIn_exceptionVec_2),
    .io_cfIn_exceptionVec_4(csr_io_cfIn_exceptionVec_4),
    .io_cfIn_exceptionVec_6(csr_io_cfIn_exceptionVec_6),
    .io_cfIn_exceptionVec_12(csr_io_cfIn_exceptionVec_12),
    .io_cfIn_intrVec_0(csr_io_cfIn_intrVec_0),
    .io_cfIn_intrVec_1(csr_io_cfIn_intrVec_1),
    .io_cfIn_intrVec_2(csr_io_cfIn_intrVec_2),
    .io_cfIn_intrVec_3(csr_io_cfIn_intrVec_3),
    .io_cfIn_intrVec_4(csr_io_cfIn_intrVec_4),
    .io_cfIn_intrVec_5(csr_io_cfIn_intrVec_5),
    .io_cfIn_intrVec_6(csr_io_cfIn_intrVec_6),
    .io_cfIn_intrVec_7(csr_io_cfIn_intrVec_7),
    .io_cfIn_intrVec_8(csr_io_cfIn_intrVec_8),
    .io_cfIn_intrVec_9(csr_io_cfIn_intrVec_9),
    .io_cfIn_intrVec_10(csr_io_cfIn_intrVec_10),
    .io_cfIn_intrVec_11(csr_io_cfIn_intrVec_11),
    .io_cfIn_crossPageIPFFix(csr_io_cfIn_crossPageIPFFix),
    .io_redirect_target(csr_io_redirect_target),
    .io_redirect_valid(csr_io_redirect_valid),
    .io_instrValid(csr_io_instrValid),
    .io_intrNO(csr_io_intrNO),
    .io_imemMMU_priviledgeMode(csr_io_imemMMU_priviledgeMode),
    .io_dmemMMU_priviledgeMode(csr_io_dmemMMU_priviledgeMode),
    .io_dmemMMU_status_sum(csr_io_dmemMMU_status_sum),
    .io_dmemMMU_status_mxr(csr_io_dmemMMU_status_mxr),
    .io_dmemMMU_loadPF(csr_io_dmemMMU_loadPF),
    .io_dmemMMU_storePF(csr_io_dmemMMU_storePF),
    .io_dmemMMU_addr(csr_io_dmemMMU_addr),
    .io_wenFix(csr_io_wenFix),
    ._T_4181_0(csr__T_4181_0),
    .perfCntCondMloadInstr(csr_perfCntCondMloadInstr),
    ._T_4184_0(csr__T_4184_0),
    .perfCntCondMlsuInstr(csr_perfCntCondMlsuInstr),
    .set_lr(csr_set_lr),
    .perfCntCondMrawStall(csr_perfCntCondMrawStall),
    .Custom4(csr_Custom4),
    .Custom7(csr_Custom7),
    ._T_4185_0(csr__T_4185_0),
    .MbpRRight(csr_MbpRRight),
    .perfCnts_2_0(csr_perfCnts_2_0),
    .satp_0(csr_satp_0),
    ._T_4178_0(csr__T_4178_0),
    .Custom6(csr_Custom6),
    .perfCntCondMinstret(csr_perfCntCondMinstret),
    .MbpBRight(csr_MbpBRight),
    .perfCntCondMexuBusy(csr_perfCntCondMexuBusy),
    .perfCntCondMmduInstr(csr_perfCntCondMmduInstr),
    .mtip_0(csr_mtip_0),
    .Custom3(csr_Custom3),
    .DISPLAY_ENABLE(csr_DISPLAY_ENABLE),
    .MbpBWrong(csr_MbpBWrong),
    .MbpRWrong(csr_MbpRWrong),
    .meip_0(csr_meip_0),
    .perfCntCondISUIssue(csr_perfCntCondISUIssue),
    .nutcoretrap_0(csr_nutcoretrap_0),
    .MbpIRight(csr_MbpIRight),
    .perfCntCondMcsrInstr(csr_perfCntCondMcsrInstr),
    .perfCntCondMsnnInstr(csr_perfCntCondMsnnInstr),
    .perfCntCondMmulInstr(csr_perfCntCondMmulInstr),
    .LSUADDR(csr_LSUADDR),
    .Custom5(csr_Custom5),
    .MbpJRight(csr_MbpJRight),
    .perfCntCondMbruInstr(csr_perfCntCondMbruInstr),
    .intrVec_0(csr_intrVec_0),
    .perfCntCondMaluInstr(csr_perfCntCondMaluInstr),
    .Custom8(csr_Custom8),
    .perfCntCondMloadStall(csr_perfCntCondMloadStall),
    .Custom2(csr_Custom2),
    .msip_0(csr_msip_0),
    .MbpIWrong(csr_MbpIWrong),
    .set_lr_addr(csr_set_lr_addr),
    .perfCntCondMimemStall(csr_perfCntCondMimemStall),
    .perfCntCondMstoreStall(csr_perfCntCondMstoreStall),
    ._T_4183_0(csr__T_4183_0),
    ._T_4182_0(csr__T_4182_0),
    .perfCnts_0_0(csr_perfCnts_0_0),
    .perfCntCondMifuFlush(csr_perfCntCondMifuFlush),
    ._T_4179_0(csr__T_4179_0),
    .perfCntCondMmmioInstr(csr_perfCntCondMmmioInstr),
    .perfCntCondMultiCommit(csr_perfCntCondMultiCommit),
    .Custom1(csr_Custom1),
    .MbpJWrong(csr_MbpJWrong),
    .set_lr_val(csr_set_lr_val),
    .lrAddr_0(csr_lrAddr_0)
  );
  MOU mou ( // @[EXU.scala 81:19]
    .clock(mou_clock),
    .reset(mou_reset),
    .io_in_valid(mou_io_in_valid),
    .io_in_bits_func(mou_io_in_bits_func),
    .io_cfIn_pc(mou_io_cfIn_pc),
    .io_redirect_target(mou_io_redirect_target),
    .io_redirect_valid(mou_io_redirect_valid),
    .flushICache_0(mou_flushICache_0),
    .DISPLAY_ENABLE(mou_DISPLAY_ENABLE),
    .flushTLB_0(mou_flushTLB_0)
  );
  SNN snn ( // @[EXU.scala 87:19]
    .clock(snn_clock),
    .reset(snn_reset),
    .io_in_valid(snn_io_in_valid),
    .io_in_bits_src1(snn_io_in_bits_src1),
    .io_in_bits_src2(snn_io_in_bits_src2),
    .io_in_bits_func(snn_io_in_bits_func),
    .io_out_ready(snn_io_out_ready),
    .io_out_valid(snn_io_out_valid),
    .io_out_bits(snn_io_out_bits),
    .io_imm(snn_io_imm),
    .io_srf_0(snn_io_srf_0),
    .io_srf_1(snn_io_srf_1),
    .io_srf_2(snn_io_srf_2),
    .io_srf_3(snn_io_srf_3),
    .io_srfAddrGen(snn_io_srfAddrGen),
    .io_wen(snn_io_wen)
  );
  Monitor Monitor ( // @[EXU.scala 144:21]
    .clk(Monitor_clk),
    .reset(Monitor_reset),
    .isNutCoreTrap(Monitor_isNutCoreTrap),
    .trapCode(Monitor_trapCode),
    .trapPC(Monitor_trapPC),
    .cycleCnt(Monitor_cycleCnt),
    .instrCnt(Monitor_instrCnt)
  );
  assign io__in_ready = _T_79 | io__out_valid; // @[EXU.scala 124:15]
  assign io__out_valid = io__in_valid & _T_77; // @[EXU.scala 111:16]
  assign io__out_bits_decode_cf_instr = io__in_bits_cf_instr; // @[EXU.scala 102:31]
  assign io__out_bits_decode_cf_pc = io__in_bits_cf_pc; // @[EXU.scala 101:28]
  assign io__out_bits_decode_cf_redirect_target = mou_io_redirect_valid ? mou_io_redirect_target : _T_48_target; // @[EXU.scala 103:34]
  assign io__out_bits_decode_cf_redirect_valid = mou_io_redirect_valid ? mou_io_redirect_valid : _T_48_valid; // @[EXU.scala 103:34]
  assign io__out_bits_decode_ctrl_fuType = io__in_bits_ctrl_fuType; // @[EXU.scala 97:14]
  assign io__out_bits_decode_ctrl_rfWen = _T_42 & _T_44; // @[EXU.scala 95:13]
  assign io__out_bits_decode_ctrl_rfDest = io__in_bits_ctrl_rfDest; // @[EXU.scala 96:14]
  assign io__out_bits_decode_ctrl_srfWen = snn_io_wen & _T_46; // @[EXU.scala 98:14]
  assign io__out_bits_decode_ctrl_srfDest = snn_io_srfAddrGen; // @[EXU.scala 99:15]
  assign io__out_bits_isMMIO = lsu_io__isMMIO | _T_31; // @[EXU.scala 58:22]
  assign io__out_bits_intrNO = csr_io_intrNO; // @[EXU.scala 74:22]
  assign io__out_bits_commits_0 = alu_io_out_bits; // @[EXU.scala 117:35]
  assign io__out_bits_commits_1 = lsu_io__out_bits; // @[EXU.scala 118:35]
  assign io__out_bits_commits_2 = mdu_io_out_bits; // @[EXU.scala 120:35]
  assign io__out_bits_commits_3 = csr_io_out_bits; // @[EXU.scala 119:35]
  assign io__out_bits_commits_5 = snn_io_out_bits; // @[EXU.scala 122:35]
  assign io__dmem_req_valid = lsu_io__dmem_req_valid; // @[EXU.scala 59:11]
  assign io__dmem_req_bits_addr = lsu_io__dmem_req_bits_addr; // @[EXU.scala 59:11]
  assign io__dmem_req_bits_size = lsu_io__dmem_req_bits_size; // @[EXU.scala 59:11]
  assign io__dmem_req_bits_cmd = lsu_io__dmem_req_bits_cmd; // @[EXU.scala 59:11]
  assign io__dmem_req_bits_wmask = lsu_io__dmem_req_bits_wmask; // @[EXU.scala 59:11]
  assign io__dmem_req_bits_wdata = lsu_io__dmem_req_bits_wdata; // @[EXU.scala 59:11]
  assign io__forward_valid = io__in_valid; // @[EXU.scala 126:20]
  assign io__forward_wb_rfWen = io__in_bits_ctrl_rfWen; // @[EXU.scala 127:23]
  assign io__forward_wb_rfDest = io__in_bits_ctrl_rfDest; // @[EXU.scala 129:24]
  assign io__forward_wb_rfData = _T_82 ? alu_io_out_bits : lsu_io__out_bits; // @[EXU.scala 131:24]
  assign io__forward_wb_srfDest = snn_io_srfAddrGen; // @[EXU.scala 130:25]
  assign io__forward_wb_srfData = snn_io_out_bits; // @[EXU.scala 132:25]
  assign io__forward_fuType = io__in_bits_ctrl_fuType; // @[EXU.scala 133:21]
  assign io__memMMU_imem_priviledgeMode = csr_io_imemMMU_priviledgeMode; // @[EXU.scala 78:18]
  assign io__memMMU_dmem_priviledgeMode = csr_io_dmemMMU_priviledgeMode; // @[EXU.scala 79:18]
  assign io__memMMU_dmem_status_sum = csr_io_dmemMMU_status_sum; // @[EXU.scala 79:18]
  assign io__memMMU_dmem_status_mxr = csr_io_dmemMMU_status_mxr; // @[EXU.scala 79:18]
  assign _T_4181 = csr__T_4181_0;
  assign _T_4184 = csr__T_4184_0;
  assign flushICache = mou_flushICache_0;
  assign _T_4185 = csr__T_4185_0;
  assign satp = csr_satp_0;
  assign _T_243_valid = alu__T_243_0_valid;
  assign _T_243_pc = alu__T_243_0_pc;
  assign _T_243_isMissPredict = alu__T_243_0_isMissPredict;
  assign _T_243_actualTarget = alu__T_243_0_actualTarget;
  assign _T_243_actualTaken = alu__T_243_0_actualTaken;
  assign _T_243_fuOpType = alu__T_243_0_fuOpType;
  assign _T_243_btbType = alu__T_243_0_btbType;
  assign _T_243_isRVC = alu__T_243_0_isRVC;
  assign _T_4178 = csr__T_4178_0;
  assign amoReq = lsu_amoReq_0;
  assign intrVec = csr_intrVec_0;
  assign _T_4183 = csr__T_4183_0;
  assign _T_4182 = csr__T_4182_0;
  assign flushTLB = mou_flushTLB_0;
  assign _T_4179 = csr__T_4179_0;
  assign alu_clock = clock;
  assign alu_reset = reset;
  assign alu_io_in_valid = _T_1 & _T_2; // @[ALU.scala 79:16]
  assign alu_io_in_bits_src1 = io__in_bits_data_src1; // @[ALU.scala 80:15]
  assign alu_io_in_bits_src2 = io__in_bits_data_src2; // @[ALU.scala 81:15]
  assign alu_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[ALU.scala 82:15]
  assign alu_io_out_ready = 1'h1; // @[EXU.scala 49:20]
  assign alu_io_cfIn_instr = io__in_bits_cf_instr; // @[EXU.scala 47:15]
  assign alu_io_cfIn_pc = io__in_bits_cf_pc; // @[EXU.scala 47:15]
  assign alu_io_cfIn_pnpc = io__in_bits_cf_pnpc; // @[EXU.scala 47:15]
  assign alu_io_cfIn_brIdx = io__in_bits_cf_brIdx; // @[EXU.scala 47:15]
  assign alu_io_offset = io__in_bits_data_imm; // @[EXU.scala 48:17]
  assign alu_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign lsu_clock = clock;
  assign lsu_reset = reset;
  assign lsu_io__in_valid = _T_5 & _T_2; // @[UnpipelinedLSU.scala 40:16]
  assign lsu_io__in_bits_src1 = io__in_bits_data_src1; // @[UnpipelinedLSU.scala 41:15]
  assign lsu_io__in_bits_src2 = io__in_bits_data_imm; // @[UnpipelinedLSU.scala 42:15]
  assign lsu_io__in_bits_func = io__in_bits_ctrl_fuOpType; // @[UnpipelinedLSU.scala 43:15]
  assign lsu_io__out_ready = 1'h1; // @[EXU.scala 60:20]
  assign lsu_io__wdata = io__in_bits_data_src2; // @[EXU.scala 56:16]
  assign lsu_io__instr = io__in_bits_cf_instr[31:0]; // @[EXU.scala 57:16]
  assign lsu_io__dmem_req_ready = io__dmem_req_ready; // @[EXU.scala 59:11]
  assign lsu_io__dmem_resp_valid = io__dmem_resp_valid; // @[EXU.scala 59:11]
  assign lsu_io__dmem_resp_bits_rdata = io__dmem_resp_bits_rdata; // @[EXU.scala 59:11]
  assign lsu_DTLBPF = _T_38_0;
  assign lsu_lsuMMIO_0 = mmio;
  assign lsu_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign lsu_DTLBENABLE = vmEnable;
  assign lsu_DTLBFINISH = _T_37_1;
  assign lsu_lr_addr = csr_lrAddr_0;
  assign mdu_clock = clock;
  assign mdu_reset = reset;
  assign mdu_io_in_valid = _T_9 & _T_2; // @[MDU.scala 140:16]
  assign mdu_io_in_bits_src1 = io__in_bits_data_src1; // @[MDU.scala 141:15]
  assign mdu_io_in_bits_src2 = io__in_bits_data_src2; // @[MDU.scala 142:15]
  assign mdu_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[MDU.scala 143:15]
  assign mdu_io_out_ready = 1'h1; // @[EXU.scala 64:20]
  assign mdu_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_in_valid = _T_13 & _T_2; // @[CSR.scala 196:16]
  assign csr_io_in_bits_src1 = io__in_bits_data_src1; // @[CSR.scala 197:15]
  assign csr_io_in_bits_src2 = io__in_bits_data_src2; // @[CSR.scala 198:15]
  assign csr_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[CSR.scala 199:15]
  assign csr_io_out_ready = 1'h1; // @[EXU.scala 76:20]
  assign csr_io_cfIn_instr = io__in_bits_cf_instr; // @[EXU.scala 69:15]
  assign csr_io_cfIn_pc = io__in_bits_cf_pc; // @[EXU.scala 69:15]
  assign csr_io_cfIn_exceptionVec_1 = io__in_bits_cf_exceptionVec_1; // @[EXU.scala 69:15]
  assign csr_io_cfIn_exceptionVec_2 = io__in_bits_cf_exceptionVec_2; // @[EXU.scala 69:15]
  assign csr_io_cfIn_exceptionVec_4 = lsu_io__loadAddrMisaligned; // @[EXU.scala 69:15 EXU.scala 70:48]
  assign csr_io_cfIn_exceptionVec_6 = lsu_io__storeAddrMisaligned; // @[EXU.scala 69:15 EXU.scala 71:49]
  assign csr_io_cfIn_exceptionVec_12 = io__in_bits_cf_exceptionVec_12; // @[EXU.scala 69:15]
  assign csr_io_cfIn_intrVec_0 = io__in_bits_cf_intrVec_0; // @[EXU.scala 69:15]
  assign csr_io_cfIn_intrVec_1 = io__in_bits_cf_intrVec_1; // @[EXU.scala 69:15]
  assign csr_io_cfIn_intrVec_2 = io__in_bits_cf_intrVec_2; // @[EXU.scala 69:15]
  assign csr_io_cfIn_intrVec_3 = io__in_bits_cf_intrVec_3; // @[EXU.scala 69:15]
  assign csr_io_cfIn_intrVec_4 = io__in_bits_cf_intrVec_4; // @[EXU.scala 69:15]
  assign csr_io_cfIn_intrVec_5 = io__in_bits_cf_intrVec_5; // @[EXU.scala 69:15]
  assign csr_io_cfIn_intrVec_6 = io__in_bits_cf_intrVec_6; // @[EXU.scala 69:15]
  assign csr_io_cfIn_intrVec_7 = io__in_bits_cf_intrVec_7; // @[EXU.scala 69:15]
  assign csr_io_cfIn_intrVec_8 = io__in_bits_cf_intrVec_8; // @[EXU.scala 69:15]
  assign csr_io_cfIn_intrVec_9 = io__in_bits_cf_intrVec_9; // @[EXU.scala 69:15]
  assign csr_io_cfIn_intrVec_10 = io__in_bits_cf_intrVec_10; // @[EXU.scala 69:15]
  assign csr_io_cfIn_intrVec_11 = io__in_bits_cf_intrVec_11; // @[EXU.scala 69:15]
  assign csr_io_cfIn_crossPageIPFFix = io__in_bits_cf_crossPageIPFFix; // @[EXU.scala 69:15]
  assign csr_io_instrValid = io__in_valid & _T_2; // @[EXU.scala 72:21]
  assign csr_io_dmemMMU_loadPF = io__memMMU_dmem_loadPF; // @[EXU.scala 79:18]
  assign csr_io_dmemMMU_storePF = io__memMMU_dmem_storePF; // @[EXU.scala 79:18]
  assign csr_io_dmemMMU_addr = io__memMMU_dmem_addr; // @[EXU.scala 79:18]
  assign csr_perfCntCondMloadInstr = lsu__T_250;
  assign csr_perfCntCondMlsuInstr = _T_89;
  assign csr_set_lr = lsu_setLr_0;
  assign csr_perfCntCondMrawStall = _T_183;
  assign csr_Custom4 = alu__T_272_0;
  assign csr_Custom7 = alu__T_288_0;
  assign csr_MbpRRight = alu__T_308_0;
  assign csr_Custom6 = alu__T_283_0;
  assign csr_perfCntCondMinstret = io_in_valid;
  assign csr_MbpBRight = alu__T_249_0;
  assign csr_perfCntCondMexuBusy = _T_186;
  assign csr_perfCntCondMmduInstr = _T_90;
  assign csr_mtip_0 = io_extra_mtip;
  assign csr_Custom3 = alu__T_266_0;
  assign csr_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign csr_MbpBWrong = alu__T_250_1;
  assign csr_MbpRWrong = alu__T_310_0;
  assign csr_meip_0 = io_extra_meip_0;
  assign csr_perfCntCondISUIssue = _T_187;
  assign csr_nutcoretrap_0 = _T_95;
  assign csr_MbpIRight = alu__T_304_0;
  assign csr_perfCntCondMcsrInstr = _T_92;
  assign csr_perfCntCondMsnnInstr = _T_91;
  assign csr_perfCntCondMmulInstr = mdu__T_87_0;
  assign csr_LSUADDR = lsu_io_in_bits_src1;
  assign csr_Custom5 = alu__T_277_0;
  assign csr_MbpJRight = alu__T_298_0;
  assign csr_perfCntCondMbruInstr = _T_88;
  assign csr_perfCntCondMaluInstr = _T_86;
  assign csr_Custom8 = alu__T_294_0;
  assign csr_perfCntCondMloadStall = lsu__T_258;
  assign csr_Custom2 = alu__T_261_0;
  assign csr_msip_0 = io_extra_msip;
  assign csr_MbpIWrong = alu__T_306_0;
  assign csr_set_lr_addr = lsu_setLrAddr_0;
  assign csr_perfCntCondMimemStall = _T_65_0;
  assign csr_perfCntCondMstoreStall = lsu__T_262;
  assign csr_perfCntCondMifuFlush = _T_66_0;
  assign csr_perfCntCondMmmioInstr = lsu_io_isMMIO;
  assign csr_perfCntCondMultiCommit = falseWire_1;
  assign csr_Custom1 = alu__T_255_0;
  assign csr_MbpJWrong = alu__T_302_0;
  assign csr_set_lr_val = lsu_setLrVal_0;
  assign mou_clock = clock;
  assign mou_reset = reset;
  assign mou_io_in_valid = _T_17 & _T_2; // @[MOU.scala 42:16]
  assign mou_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[MOU.scala 45:15]
  assign mou_io_cfIn_pc = io__in_bits_cf_pc; // @[EXU.scala 84:15]
  assign mou_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign snn_clock = clock;
  assign snn_reset = reset;
  assign snn_io_in_valid = _T_21 & _T_2; // @[SNN.scala 75:20]
  assign snn_io_in_bits_src1 = io__in_bits_data_src1; // @[SNN.scala 76:19]
  assign snn_io_in_bits_src2 = io__in_bits_data_src2; // @[SNN.scala 77:19]
  assign snn_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[SNN.scala 78:19]
  assign snn_io_out_ready = 1'h1; // @[EXU.scala 90:20]
  assign snn_io_imm = io__in_bits_data_imm; // @[EXU.scala 89:14]
  assign snn_io_srf_0 = io__in_bits_data_srf_0; // @[EXU.scala 91:15]
  assign snn_io_srf_1 = io__in_bits_data_srf_1; // @[EXU.scala 91:15]
  assign snn_io_srf_2 = io__in_bits_data_srf_2; // @[EXU.scala 91:15]
  assign snn_io_srf_3 = io__in_bits_data_srf_3; // @[EXU.scala 91:15]
  assign Monitor_clk = clock; // @[EXU.scala 148:16]
  assign Monitor_reset = reset; // @[EXU.scala 149:18]
  assign Monitor_isNutCoreTrap = _T_95; // @[EXU.scala 150:26]
  assign Monitor_trapCode = io__in_bits_data_src1[31:0]; // @[EXU.scala 151:21]
  assign Monitor_trapPC = {{25'd0}, io__in_bits_cf_pc}; // @[EXU.scala 152:19]
  assign Monitor_cycleCnt = csr_perfCnts_0_0; // @[EXU.scala 153:21]
  assign Monitor_instrCnt = csr_perfCnts_2_0; // @[EXU.scala 154:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  _T_52 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  _T_63 = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_52 <= 64'h0;
    end else begin
      _T_52 <= _T_54;
    end
    if (reset) begin
      _T_63 <= 64'h0;
    end else begin
      _T_63 <= _T_65;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_56 & _T_58) begin
          $fwrite(32'h80000002,"[%d] EXU: ",_T_52); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_56 & _T_58) begin
          $fwrite(32'h80000002,"[REDIRECT] mou %x csr %x alu %x \n",mou_io_redirect_valid,csr_io_redirect_valid,alu_io_redirect_valid); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_56 & _T_58) begin
          $fwrite(32'h80000002,"[%d] EXU: ",_T_63); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_56 & _T_58) begin
          $fwrite(32'h80000002,"[REDIRECT] flush: %d mou %x csr %x alu %x\n",io__flush,mou_io_redirect_target,csr_io_redirect_target,alu_io_redirect_target); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module WBU(
  input         clock,
  input         reset,
  input         io__in_valid,
  input  [63:0] io__in_bits_decode_cf_instr,
  input  [38:0] io__in_bits_decode_cf_pc,
  input  [38:0] io__in_bits_decode_cf_redirect_target,
  input         io__in_bits_decode_cf_redirect_valid,
  input  [2:0]  io__in_bits_decode_ctrl_fuType,
  input         io__in_bits_decode_ctrl_rfWen,
  input  [4:0]  io__in_bits_decode_ctrl_rfDest,
  input         io__in_bits_decode_ctrl_srfWen,
  input  [2:0]  io__in_bits_decode_ctrl_srfDest,
  input         io__in_bits_isMMIO,
  input  [63:0] io__in_bits_intrNO,
  input  [63:0] io__in_bits_commits_0,
  input  [63:0] io__in_bits_commits_1,
  input  [63:0] io__in_bits_commits_2,
  input  [63:0] io__in_bits_commits_3,
  input  [63:0] io__in_bits_commits_5,
  output        io__wb_rfWen,
  output [4:0]  io__wb_rfDest,
  output [63:0] io__wb_rfData,
  output        io__wb_srfWen,
  output [2:0]  io__wb_srfDest,
  output [63:0] io__wb_srfData,
  output [38:0] io__redirect_target,
  output        io__redirect_valid,
  output        falseWire_0,
  output        falseWire_1,
  output        io_in_valid,
  output        _T_36_0,
  output [63:0] _T_32_0,
  input         DISPLAY_ENABLE,
  output [63:0] _T_31_0,
  output [63:0] _T_37_0,
  output        _T_26_0,
  output        _T_33_0,
  output        falseWire_2
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] _GEN_1 = 3'h1 == io__in_bits_decode_ctrl_fuType ? io__in_bits_commits_1 : io__in_bits_commits_0; // @[WBU.scala 33:16]
  wire [63:0] _GEN_2 = 3'h2 == io__in_bits_decode_ctrl_fuType ? io__in_bits_commits_2 : _GEN_1; // @[WBU.scala 33:16]
  wire [63:0] _GEN_3 = 3'h3 == io__in_bits_decode_ctrl_fuType ? io__in_bits_commits_3 : _GEN_2; // @[WBU.scala 33:16]
  wire [63:0] _GEN_4 = 3'h4 == io__in_bits_decode_ctrl_fuType ? 64'h0 : _GEN_3; // @[WBU.scala 33:16]
  wire  _T_1 = io__in_bits_decode_ctrl_srfWen & io__in_valid; // @[WBU.scala 34:49]
  wire  _T_2 = io__in_bits_decode_ctrl_srfDest != 3'h0; // @[WBU.scala 34:99]
  wire  _T_8 = 1'h0; // @[WBU.scala 43:38]
  wire  _T_10 = ~reset; // @[WBU.scala 44:11]
  reg [63:0] _T_17; // @[GTimer.scala 24:20]
  wire [63:0] _T_19 = _T_17 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_21 = io__in_valid & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  reg  _T_26; // @[WBU.scala 57:34]
  wire [24:0] _T_29 = io__in_bits_decode_cf_pc[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  reg [63:0] _T_31; // @[WBU.scala 59:34]
  reg [63:0] _T_32; // @[WBU.scala 60:34]
  reg  _T_33; // @[WBU.scala 61:34]
  reg  _T_36; // @[WBU.scala 62:34]
  reg [63:0] _T_37; // @[WBU.scala 64:34]
  wire  falseWire = 1'h0;
  assign io__wb_rfWen = io__in_bits_decode_ctrl_rfWen & io__in_valid; // @[WBU.scala 31:15]
  assign io__wb_rfDest = io__in_bits_decode_ctrl_rfDest; // @[WBU.scala 32:16]
  assign io__wb_rfData = 3'h5 == io__in_bits_decode_ctrl_fuType ? io__in_bits_commits_5 : _GEN_4; // @[WBU.scala 33:16]
  assign io__wb_srfWen = _T_1 & _T_2; // @[WBU.scala 34:16]
  assign io__wb_srfDest = io__in_bits_decode_ctrl_srfDest; // @[WBU.scala 35:17]
  assign io__wb_srfData = _T_1 ? io__in_bits_commits_5 : 64'h0; // @[WBU.scala 36:17]
  assign io__redirect_target = io__in_bits_decode_cf_redirect_target; // @[WBU.scala 40:15]
  assign io__redirect_valid = io__in_bits_decode_cf_redirect_valid & io__in_valid; // @[WBU.scala 40:15 WBU.scala 41:21]
  assign falseWire_0 = _T_8;
  assign falseWire_1 = _T_8;
  assign io_in_valid = io__in_valid;
  assign _T_36_0 = _T_36;
  assign _T_32_0 = _T_32;
  assign _T_31_0 = _T_31;
  assign _T_37_0 = _T_37;
  assign _T_26_0 = _T_26;
  assign _T_33_0 = _T_33;
  assign falseWire_2 = _T_8;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  _T_17 = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  _T_31 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  _T_32 = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  _T_33 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _T_36 = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  _T_37 = _RAND_6[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_17 <= 64'h0;
    end else begin
      _T_17 <= _T_19;
    end
    _T_26 <= io__in_valid;
    _T_31 <= {_T_29,io__in_bits_decode_cf_pc};
    _T_32 <= io__in_bits_decode_cf_instr;
    _T_33 <= io__in_bits_isMMIO;
    _T_36 <= io__in_bits_decode_cf_instr[1:0] != 2'h3;
    _T_37 <= io__in_bits_intrNO;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_21 & _T_10) begin
          $fwrite(32'h80000002,"[%d] WBU: ",_T_17); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_21 & _T_10) begin
          $fwrite(32'h80000002,"[COMMIT] pc = 0x%x inst %x wen %x wdst %x wdata %x mmio %x intrNO %x\n",io__in_bits_decode_cf_pc,io__in_bits_decode_cf_instr,io__wb_rfWen,io__wb_rfDest,io__wb_rfData,io__in_bits_isMMIO,io__in_bits_intrNO); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Backend_inorder(
  input         clock,
  input         reset,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [63:0] io_in_0_bits_cf_instr,
  input  [38:0] io_in_0_bits_cf_pc,
  input  [38:0] io_in_0_bits_cf_pnpc,
  input         io_in_0_bits_cf_exceptionVec_1,
  input         io_in_0_bits_cf_exceptionVec_2,
  input         io_in_0_bits_cf_exceptionVec_12,
  input         io_in_0_bits_cf_intrVec_0,
  input         io_in_0_bits_cf_intrVec_1,
  input         io_in_0_bits_cf_intrVec_2,
  input         io_in_0_bits_cf_intrVec_3,
  input         io_in_0_bits_cf_intrVec_4,
  input         io_in_0_bits_cf_intrVec_5,
  input         io_in_0_bits_cf_intrVec_6,
  input         io_in_0_bits_cf_intrVec_7,
  input         io_in_0_bits_cf_intrVec_8,
  input         io_in_0_bits_cf_intrVec_9,
  input         io_in_0_bits_cf_intrVec_10,
  input         io_in_0_bits_cf_intrVec_11,
  input  [3:0]  io_in_0_bits_cf_brIdx,
  input         io_in_0_bits_cf_crossPageIPFFix,
  input  [1:0]  io_in_0_bits_ctrl_src1Type,
  input  [1:0]  io_in_0_bits_ctrl_src2Type,
  input  [2:0]  io_in_0_bits_ctrl_fuType,
  input  [6:0]  io_in_0_bits_ctrl_fuOpType,
  input  [4:0]  io_in_0_bits_ctrl_rfSrc1,
  input  [4:0]  io_in_0_bits_ctrl_rfSrc2,
  input         io_in_0_bits_ctrl_rfWen,
  input  [4:0]  io_in_0_bits_ctrl_rfDest,
  input         io_in_0_bits_ctrl_isNutCoreTrap,
  input  [63:0] io_in_0_bits_data_imm,
  input  [1:0]  io_flush,
  input         io_dmem_req_ready,
  output        io_dmem_req_valid,
  output [38:0] io_dmem_req_bits_addr,
  output [2:0]  io_dmem_req_bits_size,
  output [3:0]  io_dmem_req_bits_cmd,
  output [7:0]  io_dmem_req_bits_wmask,
  output [63:0] io_dmem_req_bits_wdata,
  input         io_dmem_resp_valid,
  input  [63:0] io_dmem_resp_bits_rdata,
  output [1:0]  io_memMMU_imem_priviledgeMode,
  output [1:0]  io_memMMU_dmem_priviledgeMode,
  output        io_memMMU_dmem_status_sum,
  output        io_memMMU_dmem_status_mxr,
  input         io_memMMU_dmem_loadPF,
  input         io_memMMU_dmem_storePF,
  input  [38:0] io_memMMU_dmem_addr,
  output [38:0] io_redirect_target,
  output        io_redirect_valid,
  output [63:0] _T_4181,
  output [63:0] _T_4184,
  input         _T_38,
  output        flushICache,
  output [63:0] _T_4185,
  output        falseWire,
  output [63:0] satp,
  output        _T_243_valid,
  output [38:0] _T_243_pc,
  output        _T_243_isMissPredict,
  output [38:0] _T_243_actualTarget,
  output        _T_243_actualTaken,
  output [6:0]  _T_243_fuOpType,
  output [1:0]  _T_243_btbType,
  output        _T_243_isRVC,
  output        falseWire_0,
  output [1:0]  _T_4178,
  output [63:0] _T_284_0,
  output [63:0] _T_284_1,
  output [63:0] _T_284_2,
  output [63:0] _T_284_3,
  output [63:0] _T_284_4,
  output [63:0] _T_284_5,
  output [63:0] _T_284_6,
  output [63:0] _T_284_7,
  output [63:0] _T_284_8,
  output [63:0] _T_284_9,
  output [63:0] _T_284_10,
  output [63:0] _T_284_11,
  output [63:0] _T_284_12,
  output [63:0] _T_284_13,
  output [63:0] _T_284_14,
  output [63:0] _T_284_15,
  output [63:0] _T_284_16,
  output [63:0] _T_284_17,
  output [63:0] _T_284_18,
  output [63:0] _T_284_19,
  output [63:0] _T_284_20,
  output [63:0] _T_284_21,
  output [63:0] _T_284_22,
  output [63:0] _T_284_23,
  output [63:0] _T_284_24,
  output [63:0] _T_284_25,
  output [63:0] _T_284_26,
  output [63:0] _T_284_27,
  output [63:0] _T_284_28,
  output [63:0] _T_284_29,
  output [63:0] _T_284_30,
  output [63:0] _T_284_31,
  input         mmio,
  output        _T_36,
  input         io_extra_mtip,
  output        amoReq,
  output [63:0] _T_32,
  input         _T_13,
  input         io_extra_meip_0,
  input         vmEnable,
  output [63:0] _T_31,
  output [63:0] _T_37,
  output        _T_26,
  output [11:0] intrVec,
  input         _T_37_0,
  input         io_extra_msip,
  input         _T_65,
  output [63:0] _T_4183,
  output [63:0] _T_4182,
  output        flushTLB,
  output        _T_33,
  input         _T_66,
  output [63:0] _T_4179
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
`endif // RANDOMIZE_REG_INIT
  wire  isu_clock; // @[Backend.scala 676:20]
  wire  isu_reset; // @[Backend.scala 676:20]
  wire  isu_io_in_0_ready; // @[Backend.scala 676:20]
  wire  isu_io_in_0_valid; // @[Backend.scala 676:20]
  wire [63:0] isu_io_in_0_bits_cf_instr; // @[Backend.scala 676:20]
  wire [38:0] isu_io_in_0_bits_cf_pc; // @[Backend.scala 676:20]
  wire [38:0] isu_io_in_0_bits_cf_pnpc; // @[Backend.scala 676:20]
  wire  isu_io_in_0_bits_cf_exceptionVec_1; // @[Backend.scala 676:20]
  wire  isu_io_in_0_bits_cf_exceptionVec_2; // @[Backend.scala 676:20]
  wire  isu_io_in_0_bits_cf_exceptionVec_12; // @[Backend.scala 676:20]
  wire  isu_io_in_0_bits_cf_intrVec_0; // @[Backend.scala 676:20]
  wire  isu_io_in_0_bits_cf_intrVec_1; // @[Backend.scala 676:20]
  wire  isu_io_in_0_bits_cf_intrVec_2; // @[Backend.scala 676:20]
  wire  isu_io_in_0_bits_cf_intrVec_3; // @[Backend.scala 676:20]
  wire  isu_io_in_0_bits_cf_intrVec_4; // @[Backend.scala 676:20]
  wire  isu_io_in_0_bits_cf_intrVec_5; // @[Backend.scala 676:20]
  wire  isu_io_in_0_bits_cf_intrVec_6; // @[Backend.scala 676:20]
  wire  isu_io_in_0_bits_cf_intrVec_7; // @[Backend.scala 676:20]
  wire  isu_io_in_0_bits_cf_intrVec_8; // @[Backend.scala 676:20]
  wire  isu_io_in_0_bits_cf_intrVec_9; // @[Backend.scala 676:20]
  wire  isu_io_in_0_bits_cf_intrVec_10; // @[Backend.scala 676:20]
  wire  isu_io_in_0_bits_cf_intrVec_11; // @[Backend.scala 676:20]
  wire [3:0] isu_io_in_0_bits_cf_brIdx; // @[Backend.scala 676:20]
  wire  isu_io_in_0_bits_cf_crossPageIPFFix; // @[Backend.scala 676:20]
  wire [1:0] isu_io_in_0_bits_ctrl_src1Type; // @[Backend.scala 676:20]
  wire [1:0] isu_io_in_0_bits_ctrl_src2Type; // @[Backend.scala 676:20]
  wire [2:0] isu_io_in_0_bits_ctrl_fuType; // @[Backend.scala 676:20]
  wire [6:0] isu_io_in_0_bits_ctrl_fuOpType; // @[Backend.scala 676:20]
  wire [4:0] isu_io_in_0_bits_ctrl_rfSrc1; // @[Backend.scala 676:20]
  wire [4:0] isu_io_in_0_bits_ctrl_rfSrc2; // @[Backend.scala 676:20]
  wire  isu_io_in_0_bits_ctrl_rfWen; // @[Backend.scala 676:20]
  wire [4:0] isu_io_in_0_bits_ctrl_rfDest; // @[Backend.scala 676:20]
  wire  isu_io_in_0_bits_ctrl_isNutCoreTrap; // @[Backend.scala 676:20]
  wire [63:0] isu_io_in_0_bits_data_imm; // @[Backend.scala 676:20]
  wire  isu_io_out_ready; // @[Backend.scala 676:20]
  wire  isu_io_out_valid; // @[Backend.scala 676:20]
  wire [63:0] isu_io_out_bits_cf_instr; // @[Backend.scala 676:20]
  wire [38:0] isu_io_out_bits_cf_pc; // @[Backend.scala 676:20]
  wire [38:0] isu_io_out_bits_cf_pnpc; // @[Backend.scala 676:20]
  wire  isu_io_out_bits_cf_exceptionVec_1; // @[Backend.scala 676:20]
  wire  isu_io_out_bits_cf_exceptionVec_2; // @[Backend.scala 676:20]
  wire  isu_io_out_bits_cf_exceptionVec_12; // @[Backend.scala 676:20]
  wire  isu_io_out_bits_cf_intrVec_0; // @[Backend.scala 676:20]
  wire  isu_io_out_bits_cf_intrVec_1; // @[Backend.scala 676:20]
  wire  isu_io_out_bits_cf_intrVec_2; // @[Backend.scala 676:20]
  wire  isu_io_out_bits_cf_intrVec_3; // @[Backend.scala 676:20]
  wire  isu_io_out_bits_cf_intrVec_4; // @[Backend.scala 676:20]
  wire  isu_io_out_bits_cf_intrVec_5; // @[Backend.scala 676:20]
  wire  isu_io_out_bits_cf_intrVec_6; // @[Backend.scala 676:20]
  wire  isu_io_out_bits_cf_intrVec_7; // @[Backend.scala 676:20]
  wire  isu_io_out_bits_cf_intrVec_8; // @[Backend.scala 676:20]
  wire  isu_io_out_bits_cf_intrVec_9; // @[Backend.scala 676:20]
  wire  isu_io_out_bits_cf_intrVec_10; // @[Backend.scala 676:20]
  wire  isu_io_out_bits_cf_intrVec_11; // @[Backend.scala 676:20]
  wire [3:0] isu_io_out_bits_cf_brIdx; // @[Backend.scala 676:20]
  wire  isu_io_out_bits_cf_crossPageIPFFix; // @[Backend.scala 676:20]
  wire [2:0] isu_io_out_bits_ctrl_fuType; // @[Backend.scala 676:20]
  wire [6:0] isu_io_out_bits_ctrl_fuOpType; // @[Backend.scala 676:20]
  wire  isu_io_out_bits_ctrl_rfWen; // @[Backend.scala 676:20]
  wire [4:0] isu_io_out_bits_ctrl_rfDest; // @[Backend.scala 676:20]
  wire  isu_io_out_bits_ctrl_isNutCoreTrap; // @[Backend.scala 676:20]
  wire [63:0] isu_io_out_bits_data_src1; // @[Backend.scala 676:20]
  wire [63:0] isu_io_out_bits_data_src2; // @[Backend.scala 676:20]
  wire [63:0] isu_io_out_bits_data_imm; // @[Backend.scala 676:20]
  wire [63:0] isu_io_out_bits_data_srf_0; // @[Backend.scala 676:20]
  wire [63:0] isu_io_out_bits_data_srf_1; // @[Backend.scala 676:20]
  wire [63:0] isu_io_out_bits_data_srf_2; // @[Backend.scala 676:20]
  wire [63:0] isu_io_out_bits_data_srf_3; // @[Backend.scala 676:20]
  wire  isu_io_wb_rfWen; // @[Backend.scala 676:20]
  wire [4:0] isu_io_wb_rfDest; // @[Backend.scala 676:20]
  wire [63:0] isu_io_wb_rfData; // @[Backend.scala 676:20]
  wire  isu_io_wb_srfWen; // @[Backend.scala 676:20]
  wire [2:0] isu_io_wb_srfDest; // @[Backend.scala 676:20]
  wire [63:0] isu_io_wb_srfData; // @[Backend.scala 676:20]
  wire  isu_io_forward_valid; // @[Backend.scala 676:20]
  wire  isu_io_forward_wb_rfWen; // @[Backend.scala 676:20]
  wire [4:0] isu_io_forward_wb_rfDest; // @[Backend.scala 676:20]
  wire [63:0] isu_io_forward_wb_rfData; // @[Backend.scala 676:20]
  wire [2:0] isu_io_forward_wb_srfDest; // @[Backend.scala 676:20]
  wire [63:0] isu_io_forward_wb_srfData; // @[Backend.scala 676:20]
  wire [2:0] isu_io_forward_fuType; // @[Backend.scala 676:20]
  wire  isu_io_flush; // @[Backend.scala 676:20]
  wire  isu__T_183_0; // @[Backend.scala 676:20]
  wire [63:0] isu__T_284_0_0; // @[Backend.scala 676:20]
  wire [63:0] isu__T_284_0_1; // @[Backend.scala 676:20]
  wire [63:0] isu__T_284_0_2; // @[Backend.scala 676:20]
  wire [63:0] isu__T_284_0_3; // @[Backend.scala 676:20]
  wire [63:0] isu__T_284_0_4; // @[Backend.scala 676:20]
  wire [63:0] isu__T_284_0_5; // @[Backend.scala 676:20]
  wire [63:0] isu__T_284_0_6; // @[Backend.scala 676:20]
  wire [63:0] isu__T_284_0_7; // @[Backend.scala 676:20]
  wire [63:0] isu__T_284_0_8; // @[Backend.scala 676:20]
  wire [63:0] isu__T_284_0_9; // @[Backend.scala 676:20]
  wire [63:0] isu__T_284_0_10; // @[Backend.scala 676:20]
  wire [63:0] isu__T_284_0_11; // @[Backend.scala 676:20]
  wire [63:0] isu__T_284_0_12; // @[Backend.scala 676:20]
  wire [63:0] isu__T_284_0_13; // @[Backend.scala 676:20]
  wire [63:0] isu__T_284_0_14; // @[Backend.scala 676:20]
  wire [63:0] isu__T_284_0_15; // @[Backend.scala 676:20]
  wire [63:0] isu__T_284_0_16; // @[Backend.scala 676:20]
  wire [63:0] isu__T_284_0_17; // @[Backend.scala 676:20]
  wire [63:0] isu__T_284_0_18; // @[Backend.scala 676:20]
  wire [63:0] isu__T_284_0_19; // @[Backend.scala 676:20]
  wire [63:0] isu__T_284_0_20; // @[Backend.scala 676:20]
  wire [63:0] isu__T_284_0_21; // @[Backend.scala 676:20]
  wire [63:0] isu__T_284_0_22; // @[Backend.scala 676:20]
  wire [63:0] isu__T_284_0_23; // @[Backend.scala 676:20]
  wire [63:0] isu__T_284_0_24; // @[Backend.scala 676:20]
  wire [63:0] isu__T_284_0_25; // @[Backend.scala 676:20]
  wire [63:0] isu__T_284_0_26; // @[Backend.scala 676:20]
  wire [63:0] isu__T_284_0_27; // @[Backend.scala 676:20]
  wire [63:0] isu__T_284_0_28; // @[Backend.scala 676:20]
  wire [63:0] isu__T_284_0_29; // @[Backend.scala 676:20]
  wire [63:0] isu__T_284_0_30; // @[Backend.scala 676:20]
  wire [63:0] isu__T_284_0_31; // @[Backend.scala 676:20]
  wire  isu__T_186_0; // @[Backend.scala 676:20]
  wire  isu_DISPLAY_ENABLE; // @[Backend.scala 676:20]
  wire  isu__T_187_0; // @[Backend.scala 676:20]
  wire  exu_clock; // @[Backend.scala 677:20]
  wire  exu_reset; // @[Backend.scala 677:20]
  wire  exu_io__in_ready; // @[Backend.scala 677:20]
  wire  exu_io__in_valid; // @[Backend.scala 677:20]
  wire [63:0] exu_io__in_bits_cf_instr; // @[Backend.scala 677:20]
  wire [38:0] exu_io__in_bits_cf_pc; // @[Backend.scala 677:20]
  wire [38:0] exu_io__in_bits_cf_pnpc; // @[Backend.scala 677:20]
  wire  exu_io__in_bits_cf_exceptionVec_1; // @[Backend.scala 677:20]
  wire  exu_io__in_bits_cf_exceptionVec_2; // @[Backend.scala 677:20]
  wire  exu_io__in_bits_cf_exceptionVec_12; // @[Backend.scala 677:20]
  wire  exu_io__in_bits_cf_intrVec_0; // @[Backend.scala 677:20]
  wire  exu_io__in_bits_cf_intrVec_1; // @[Backend.scala 677:20]
  wire  exu_io__in_bits_cf_intrVec_2; // @[Backend.scala 677:20]
  wire  exu_io__in_bits_cf_intrVec_3; // @[Backend.scala 677:20]
  wire  exu_io__in_bits_cf_intrVec_4; // @[Backend.scala 677:20]
  wire  exu_io__in_bits_cf_intrVec_5; // @[Backend.scala 677:20]
  wire  exu_io__in_bits_cf_intrVec_6; // @[Backend.scala 677:20]
  wire  exu_io__in_bits_cf_intrVec_7; // @[Backend.scala 677:20]
  wire  exu_io__in_bits_cf_intrVec_8; // @[Backend.scala 677:20]
  wire  exu_io__in_bits_cf_intrVec_9; // @[Backend.scala 677:20]
  wire  exu_io__in_bits_cf_intrVec_10; // @[Backend.scala 677:20]
  wire  exu_io__in_bits_cf_intrVec_11; // @[Backend.scala 677:20]
  wire [3:0] exu_io__in_bits_cf_brIdx; // @[Backend.scala 677:20]
  wire  exu_io__in_bits_cf_crossPageIPFFix; // @[Backend.scala 677:20]
  wire [2:0] exu_io__in_bits_ctrl_fuType; // @[Backend.scala 677:20]
  wire [6:0] exu_io__in_bits_ctrl_fuOpType; // @[Backend.scala 677:20]
  wire  exu_io__in_bits_ctrl_rfWen; // @[Backend.scala 677:20]
  wire [4:0] exu_io__in_bits_ctrl_rfDest; // @[Backend.scala 677:20]
  wire  exu_io__in_bits_ctrl_isNutCoreTrap; // @[Backend.scala 677:20]
  wire [63:0] exu_io__in_bits_data_src1; // @[Backend.scala 677:20]
  wire [63:0] exu_io__in_bits_data_src2; // @[Backend.scala 677:20]
  wire [63:0] exu_io__in_bits_data_imm; // @[Backend.scala 677:20]
  wire [63:0] exu_io__in_bits_data_srf_0; // @[Backend.scala 677:20]
  wire [63:0] exu_io__in_bits_data_srf_1; // @[Backend.scala 677:20]
  wire [63:0] exu_io__in_bits_data_srf_2; // @[Backend.scala 677:20]
  wire [63:0] exu_io__in_bits_data_srf_3; // @[Backend.scala 677:20]
  wire  exu_io__out_ready; // @[Backend.scala 677:20]
  wire  exu_io__out_valid; // @[Backend.scala 677:20]
  wire [63:0] exu_io__out_bits_decode_cf_instr; // @[Backend.scala 677:20]
  wire [38:0] exu_io__out_bits_decode_cf_pc; // @[Backend.scala 677:20]
  wire [38:0] exu_io__out_bits_decode_cf_redirect_target; // @[Backend.scala 677:20]
  wire  exu_io__out_bits_decode_cf_redirect_valid; // @[Backend.scala 677:20]
  wire [2:0] exu_io__out_bits_decode_ctrl_fuType; // @[Backend.scala 677:20]
  wire  exu_io__out_bits_decode_ctrl_rfWen; // @[Backend.scala 677:20]
  wire [4:0] exu_io__out_bits_decode_ctrl_rfDest; // @[Backend.scala 677:20]
  wire  exu_io__out_bits_decode_ctrl_srfWen; // @[Backend.scala 677:20]
  wire [2:0] exu_io__out_bits_decode_ctrl_srfDest; // @[Backend.scala 677:20]
  wire  exu_io__out_bits_isMMIO; // @[Backend.scala 677:20]
  wire [63:0] exu_io__out_bits_intrNO; // @[Backend.scala 677:20]
  wire [63:0] exu_io__out_bits_commits_0; // @[Backend.scala 677:20]
  wire [63:0] exu_io__out_bits_commits_1; // @[Backend.scala 677:20]
  wire [63:0] exu_io__out_bits_commits_2; // @[Backend.scala 677:20]
  wire [63:0] exu_io__out_bits_commits_3; // @[Backend.scala 677:20]
  wire [63:0] exu_io__out_bits_commits_5; // @[Backend.scala 677:20]
  wire  exu_io__flush; // @[Backend.scala 677:20]
  wire  exu_io__dmem_req_ready; // @[Backend.scala 677:20]
  wire  exu_io__dmem_req_valid; // @[Backend.scala 677:20]
  wire [38:0] exu_io__dmem_req_bits_addr; // @[Backend.scala 677:20]
  wire [2:0] exu_io__dmem_req_bits_size; // @[Backend.scala 677:20]
  wire [3:0] exu_io__dmem_req_bits_cmd; // @[Backend.scala 677:20]
  wire [7:0] exu_io__dmem_req_bits_wmask; // @[Backend.scala 677:20]
  wire [63:0] exu_io__dmem_req_bits_wdata; // @[Backend.scala 677:20]
  wire  exu_io__dmem_resp_valid; // @[Backend.scala 677:20]
  wire [63:0] exu_io__dmem_resp_bits_rdata; // @[Backend.scala 677:20]
  wire  exu_io__forward_valid; // @[Backend.scala 677:20]
  wire  exu_io__forward_wb_rfWen; // @[Backend.scala 677:20]
  wire [4:0] exu_io__forward_wb_rfDest; // @[Backend.scala 677:20]
  wire [63:0] exu_io__forward_wb_rfData; // @[Backend.scala 677:20]
  wire [2:0] exu_io__forward_wb_srfDest; // @[Backend.scala 677:20]
  wire [63:0] exu_io__forward_wb_srfData; // @[Backend.scala 677:20]
  wire [2:0] exu_io__forward_fuType; // @[Backend.scala 677:20]
  wire [1:0] exu_io__memMMU_imem_priviledgeMode; // @[Backend.scala 677:20]
  wire [1:0] exu_io__memMMU_dmem_priviledgeMode; // @[Backend.scala 677:20]
  wire  exu_io__memMMU_dmem_status_sum; // @[Backend.scala 677:20]
  wire  exu_io__memMMU_dmem_status_mxr; // @[Backend.scala 677:20]
  wire  exu_io__memMMU_dmem_loadPF; // @[Backend.scala 677:20]
  wire  exu_io__memMMU_dmem_storePF; // @[Backend.scala 677:20]
  wire [38:0] exu_io__memMMU_dmem_addr; // @[Backend.scala 677:20]
  wire [63:0] exu__T_4181; // @[Backend.scala 677:20]
  wire [63:0] exu__T_4184; // @[Backend.scala 677:20]
  wire  exu__T_183; // @[Backend.scala 677:20]
  wire  exu__T_38_0; // @[Backend.scala 677:20]
  wire  exu_flushICache; // @[Backend.scala 677:20]
  wire [63:0] exu__T_4185; // @[Backend.scala 677:20]
  wire [63:0] exu_satp; // @[Backend.scala 677:20]
  wire  exu__T_243_valid; // @[Backend.scala 677:20]
  wire [38:0] exu__T_243_pc; // @[Backend.scala 677:20]
  wire  exu__T_243_isMissPredict; // @[Backend.scala 677:20]
  wire [38:0] exu__T_243_actualTarget; // @[Backend.scala 677:20]
  wire  exu__T_243_actualTaken; // @[Backend.scala 677:20]
  wire [6:0] exu__T_243_fuOpType; // @[Backend.scala 677:20]
  wire [1:0] exu__T_243_btbType; // @[Backend.scala 677:20]
  wire  exu__T_243_isRVC; // @[Backend.scala 677:20]
  wire [1:0] exu__T_4178; // @[Backend.scala 677:20]
  wire  exu_io_in_valid; // @[Backend.scala 677:20]
  wire  exu_mmio; // @[Backend.scala 677:20]
  wire  exu__T_186; // @[Backend.scala 677:20]
  wire  exu_io_extra_mtip; // @[Backend.scala 677:20]
  wire  exu_amoReq; // @[Backend.scala 677:20]
  wire  exu_DISPLAY_ENABLE; // @[Backend.scala 677:20]
  wire  exu_io_extra_meip_0; // @[Backend.scala 677:20]
  wire  exu__T_187; // @[Backend.scala 677:20]
  wire  exu_vmEnable; // @[Backend.scala 677:20]
  wire [11:0] exu_intrVec; // @[Backend.scala 677:20]
  wire  exu__T_37_1; // @[Backend.scala 677:20]
  wire  exu_io_extra_msip; // @[Backend.scala 677:20]
  wire  exu__T_65_0; // @[Backend.scala 677:20]
  wire [63:0] exu__T_4183; // @[Backend.scala 677:20]
  wire [63:0] exu__T_4182; // @[Backend.scala 677:20]
  wire  exu_flushTLB; // @[Backend.scala 677:20]
  wire  exu__T_66_0; // @[Backend.scala 677:20]
  wire [63:0] exu__T_4179; // @[Backend.scala 677:20]
  wire  exu_falseWire_1; // @[Backend.scala 677:20]
  wire  wbu_clock; // @[Backend.scala 678:20]
  wire  wbu_reset; // @[Backend.scala 678:20]
  wire  wbu_io__in_valid; // @[Backend.scala 678:20]
  wire [63:0] wbu_io__in_bits_decode_cf_instr; // @[Backend.scala 678:20]
  wire [38:0] wbu_io__in_bits_decode_cf_pc; // @[Backend.scala 678:20]
  wire [38:0] wbu_io__in_bits_decode_cf_redirect_target; // @[Backend.scala 678:20]
  wire  wbu_io__in_bits_decode_cf_redirect_valid; // @[Backend.scala 678:20]
  wire [2:0] wbu_io__in_bits_decode_ctrl_fuType; // @[Backend.scala 678:20]
  wire  wbu_io__in_bits_decode_ctrl_rfWen; // @[Backend.scala 678:20]
  wire [4:0] wbu_io__in_bits_decode_ctrl_rfDest; // @[Backend.scala 678:20]
  wire  wbu_io__in_bits_decode_ctrl_srfWen; // @[Backend.scala 678:20]
  wire [2:0] wbu_io__in_bits_decode_ctrl_srfDest; // @[Backend.scala 678:20]
  wire  wbu_io__in_bits_isMMIO; // @[Backend.scala 678:20]
  wire [63:0] wbu_io__in_bits_intrNO; // @[Backend.scala 678:20]
  wire [63:0] wbu_io__in_bits_commits_0; // @[Backend.scala 678:20]
  wire [63:0] wbu_io__in_bits_commits_1; // @[Backend.scala 678:20]
  wire [63:0] wbu_io__in_bits_commits_2; // @[Backend.scala 678:20]
  wire [63:0] wbu_io__in_bits_commits_3; // @[Backend.scala 678:20]
  wire [63:0] wbu_io__in_bits_commits_5; // @[Backend.scala 678:20]
  wire  wbu_io__wb_rfWen; // @[Backend.scala 678:20]
  wire [4:0] wbu_io__wb_rfDest; // @[Backend.scala 678:20]
  wire [63:0] wbu_io__wb_rfData; // @[Backend.scala 678:20]
  wire  wbu_io__wb_srfWen; // @[Backend.scala 678:20]
  wire [2:0] wbu_io__wb_srfDest; // @[Backend.scala 678:20]
  wire [63:0] wbu_io__wb_srfData; // @[Backend.scala 678:20]
  wire [38:0] wbu_io__redirect_target; // @[Backend.scala 678:20]
  wire  wbu_io__redirect_valid; // @[Backend.scala 678:20]
  wire  wbu_falseWire_0; // @[Backend.scala 678:20]
  wire  wbu_falseWire_1; // @[Backend.scala 678:20]
  wire  wbu_io_in_valid; // @[Backend.scala 678:20]
  wire  wbu__T_36_0; // @[Backend.scala 678:20]
  wire [63:0] wbu__T_32_0; // @[Backend.scala 678:20]
  wire  wbu_DISPLAY_ENABLE; // @[Backend.scala 678:20]
  wire [63:0] wbu__T_31_0; // @[Backend.scala 678:20]
  wire [63:0] wbu__T_37_0; // @[Backend.scala 678:20]
  wire  wbu__T_26_0; // @[Backend.scala 678:20]
  wire  wbu__T_33_0; // @[Backend.scala 678:20]
  wire  wbu_falseWire_2; // @[Backend.scala 678:20]
  wire  _T = exu_io__out_ready & exu_io__out_valid; // @[Decoupled.scala 40:37]
  reg  _T_2; // @[Pipeline.scala 24:24]
  wire  _GEN_0 = _T ? 1'h0 : _T_2; // @[Pipeline.scala 25:25]
  wire  _T_3 = isu_io_out_valid & exu_io__in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_1 = _T_3 | _GEN_0; // @[Pipeline.scala 26:38]
  reg [63:0] _T_5_cf_instr; // @[Reg.scala 15:16]
  reg [38:0] _T_5_cf_pc; // @[Reg.scala 15:16]
  reg [38:0] _T_5_cf_pnpc; // @[Reg.scala 15:16]
  reg  _T_5_cf_exceptionVec_1; // @[Reg.scala 15:16]
  reg  _T_5_cf_exceptionVec_2; // @[Reg.scala 15:16]
  reg  _T_5_cf_exceptionVec_12; // @[Reg.scala 15:16]
  reg  _T_5_cf_intrVec_0; // @[Reg.scala 15:16]
  reg  _T_5_cf_intrVec_1; // @[Reg.scala 15:16]
  reg  _T_5_cf_intrVec_2; // @[Reg.scala 15:16]
  reg  _T_5_cf_intrVec_3; // @[Reg.scala 15:16]
  reg  _T_5_cf_intrVec_4; // @[Reg.scala 15:16]
  reg  _T_5_cf_intrVec_5; // @[Reg.scala 15:16]
  reg  _T_5_cf_intrVec_6; // @[Reg.scala 15:16]
  reg  _T_5_cf_intrVec_7; // @[Reg.scala 15:16]
  reg  _T_5_cf_intrVec_8; // @[Reg.scala 15:16]
  reg  _T_5_cf_intrVec_9; // @[Reg.scala 15:16]
  reg  _T_5_cf_intrVec_10; // @[Reg.scala 15:16]
  reg  _T_5_cf_intrVec_11; // @[Reg.scala 15:16]
  reg [3:0] _T_5_cf_brIdx; // @[Reg.scala 15:16]
  reg  _T_5_cf_crossPageIPFFix; // @[Reg.scala 15:16]
  reg [2:0] _T_5_ctrl_fuType; // @[Reg.scala 15:16]
  reg [6:0] _T_5_ctrl_fuOpType; // @[Reg.scala 15:16]
  reg  _T_5_ctrl_rfWen; // @[Reg.scala 15:16]
  reg [4:0] _T_5_ctrl_rfDest; // @[Reg.scala 15:16]
  reg  _T_5_ctrl_isNutCoreTrap; // @[Reg.scala 15:16]
  reg [63:0] _T_5_data_src1; // @[Reg.scala 15:16]
  reg [63:0] _T_5_data_src2; // @[Reg.scala 15:16]
  reg [63:0] _T_5_data_imm; // @[Reg.scala 15:16]
  reg [63:0] _T_5_data_srf_0; // @[Reg.scala 15:16]
  reg [63:0] _T_5_data_srf_1; // @[Reg.scala 15:16]
  reg [63:0] _T_5_data_srf_2; // @[Reg.scala 15:16]
  reg [63:0] _T_5_data_srf_3; // @[Reg.scala 15:16]
  reg  _T_7; // @[Pipeline.scala 24:24]
  wire  _T_8 = exu_io__out_valid; // @[Pipeline.scala 26:22]
  reg [63:0] _T_10_decode_cf_instr; // @[Reg.scala 15:16]
  reg [38:0] _T_10_decode_cf_pc; // @[Reg.scala 15:16]
  reg [38:0] _T_10_decode_cf_redirect_target; // @[Reg.scala 15:16]
  reg  _T_10_decode_cf_redirect_valid; // @[Reg.scala 15:16]
  reg [2:0] _T_10_decode_ctrl_fuType; // @[Reg.scala 15:16]
  reg  _T_10_decode_ctrl_rfWen; // @[Reg.scala 15:16]
  reg [4:0] _T_10_decode_ctrl_rfDest; // @[Reg.scala 15:16]
  reg  _T_10_decode_ctrl_srfWen; // @[Reg.scala 15:16]
  reg [2:0] _T_10_decode_ctrl_srfDest; // @[Reg.scala 15:16]
  reg  _T_10_isMMIO; // @[Reg.scala 15:16]
  reg [63:0] _T_10_intrNO; // @[Reg.scala 15:16]
  reg [63:0] _T_10_commits_0; // @[Reg.scala 15:16]
  reg [63:0] _T_10_commits_1; // @[Reg.scala 15:16]
  reg [63:0] _T_10_commits_2; // @[Reg.scala 15:16]
  reg [63:0] _T_10_commits_3; // @[Reg.scala 15:16]
  reg [63:0] _T_10_commits_5; // @[Reg.scala 15:16]
  ISU isu ( // @[Backend.scala 676:20]
    .clock(isu_clock),
    .reset(isu_reset),
    .io_in_0_ready(isu_io_in_0_ready),
    .io_in_0_valid(isu_io_in_0_valid),
    .io_in_0_bits_cf_instr(isu_io_in_0_bits_cf_instr),
    .io_in_0_bits_cf_pc(isu_io_in_0_bits_cf_pc),
    .io_in_0_bits_cf_pnpc(isu_io_in_0_bits_cf_pnpc),
    .io_in_0_bits_cf_exceptionVec_1(isu_io_in_0_bits_cf_exceptionVec_1),
    .io_in_0_bits_cf_exceptionVec_2(isu_io_in_0_bits_cf_exceptionVec_2),
    .io_in_0_bits_cf_exceptionVec_12(isu_io_in_0_bits_cf_exceptionVec_12),
    .io_in_0_bits_cf_intrVec_0(isu_io_in_0_bits_cf_intrVec_0),
    .io_in_0_bits_cf_intrVec_1(isu_io_in_0_bits_cf_intrVec_1),
    .io_in_0_bits_cf_intrVec_2(isu_io_in_0_bits_cf_intrVec_2),
    .io_in_0_bits_cf_intrVec_3(isu_io_in_0_bits_cf_intrVec_3),
    .io_in_0_bits_cf_intrVec_4(isu_io_in_0_bits_cf_intrVec_4),
    .io_in_0_bits_cf_intrVec_5(isu_io_in_0_bits_cf_intrVec_5),
    .io_in_0_bits_cf_intrVec_6(isu_io_in_0_bits_cf_intrVec_6),
    .io_in_0_bits_cf_intrVec_7(isu_io_in_0_bits_cf_intrVec_7),
    .io_in_0_bits_cf_intrVec_8(isu_io_in_0_bits_cf_intrVec_8),
    .io_in_0_bits_cf_intrVec_9(isu_io_in_0_bits_cf_intrVec_9),
    .io_in_0_bits_cf_intrVec_10(isu_io_in_0_bits_cf_intrVec_10),
    .io_in_0_bits_cf_intrVec_11(isu_io_in_0_bits_cf_intrVec_11),
    .io_in_0_bits_cf_brIdx(isu_io_in_0_bits_cf_brIdx),
    .io_in_0_bits_cf_crossPageIPFFix(isu_io_in_0_bits_cf_crossPageIPFFix),
    .io_in_0_bits_ctrl_src1Type(isu_io_in_0_bits_ctrl_src1Type),
    .io_in_0_bits_ctrl_src2Type(isu_io_in_0_bits_ctrl_src2Type),
    .io_in_0_bits_ctrl_fuType(isu_io_in_0_bits_ctrl_fuType),
    .io_in_0_bits_ctrl_fuOpType(isu_io_in_0_bits_ctrl_fuOpType),
    .io_in_0_bits_ctrl_rfSrc1(isu_io_in_0_bits_ctrl_rfSrc1),
    .io_in_0_bits_ctrl_rfSrc2(isu_io_in_0_bits_ctrl_rfSrc2),
    .io_in_0_bits_ctrl_rfWen(isu_io_in_0_bits_ctrl_rfWen),
    .io_in_0_bits_ctrl_rfDest(isu_io_in_0_bits_ctrl_rfDest),
    .io_in_0_bits_ctrl_isNutCoreTrap(isu_io_in_0_bits_ctrl_isNutCoreTrap),
    .io_in_0_bits_data_imm(isu_io_in_0_bits_data_imm),
    .io_out_ready(isu_io_out_ready),
    .io_out_valid(isu_io_out_valid),
    .io_out_bits_cf_instr(isu_io_out_bits_cf_instr),
    .io_out_bits_cf_pc(isu_io_out_bits_cf_pc),
    .io_out_bits_cf_pnpc(isu_io_out_bits_cf_pnpc),
    .io_out_bits_cf_exceptionVec_1(isu_io_out_bits_cf_exceptionVec_1),
    .io_out_bits_cf_exceptionVec_2(isu_io_out_bits_cf_exceptionVec_2),
    .io_out_bits_cf_exceptionVec_12(isu_io_out_bits_cf_exceptionVec_12),
    .io_out_bits_cf_intrVec_0(isu_io_out_bits_cf_intrVec_0),
    .io_out_bits_cf_intrVec_1(isu_io_out_bits_cf_intrVec_1),
    .io_out_bits_cf_intrVec_2(isu_io_out_bits_cf_intrVec_2),
    .io_out_bits_cf_intrVec_3(isu_io_out_bits_cf_intrVec_3),
    .io_out_bits_cf_intrVec_4(isu_io_out_bits_cf_intrVec_4),
    .io_out_bits_cf_intrVec_5(isu_io_out_bits_cf_intrVec_5),
    .io_out_bits_cf_intrVec_6(isu_io_out_bits_cf_intrVec_6),
    .io_out_bits_cf_intrVec_7(isu_io_out_bits_cf_intrVec_7),
    .io_out_bits_cf_intrVec_8(isu_io_out_bits_cf_intrVec_8),
    .io_out_bits_cf_intrVec_9(isu_io_out_bits_cf_intrVec_9),
    .io_out_bits_cf_intrVec_10(isu_io_out_bits_cf_intrVec_10),
    .io_out_bits_cf_intrVec_11(isu_io_out_bits_cf_intrVec_11),
    .io_out_bits_cf_brIdx(isu_io_out_bits_cf_brIdx),
    .io_out_bits_cf_crossPageIPFFix(isu_io_out_bits_cf_crossPageIPFFix),
    .io_out_bits_ctrl_fuType(isu_io_out_bits_ctrl_fuType),
    .io_out_bits_ctrl_fuOpType(isu_io_out_bits_ctrl_fuOpType),
    .io_out_bits_ctrl_rfWen(isu_io_out_bits_ctrl_rfWen),
    .io_out_bits_ctrl_rfDest(isu_io_out_bits_ctrl_rfDest),
    .io_out_bits_ctrl_isNutCoreTrap(isu_io_out_bits_ctrl_isNutCoreTrap),
    .io_out_bits_data_src1(isu_io_out_bits_data_src1),
    .io_out_bits_data_src2(isu_io_out_bits_data_src2),
    .io_out_bits_data_imm(isu_io_out_bits_data_imm),
    .io_out_bits_data_srf_0(isu_io_out_bits_data_srf_0),
    .io_out_bits_data_srf_1(isu_io_out_bits_data_srf_1),
    .io_out_bits_data_srf_2(isu_io_out_bits_data_srf_2),
    .io_out_bits_data_srf_3(isu_io_out_bits_data_srf_3),
    .io_wb_rfWen(isu_io_wb_rfWen),
    .io_wb_rfDest(isu_io_wb_rfDest),
    .io_wb_rfData(isu_io_wb_rfData),
    .io_wb_srfWen(isu_io_wb_srfWen),
    .io_wb_srfDest(isu_io_wb_srfDest),
    .io_wb_srfData(isu_io_wb_srfData),
    .io_forward_valid(isu_io_forward_valid),
    .io_forward_wb_rfWen(isu_io_forward_wb_rfWen),
    .io_forward_wb_rfDest(isu_io_forward_wb_rfDest),
    .io_forward_wb_rfData(isu_io_forward_wb_rfData),
    .io_forward_wb_srfDest(isu_io_forward_wb_srfDest),
    .io_forward_wb_srfData(isu_io_forward_wb_srfData),
    .io_forward_fuType(isu_io_forward_fuType),
    .io_flush(isu_io_flush),
    ._T_183_0(isu__T_183_0),
    ._T_284_0_0(isu__T_284_0_0),
    ._T_284_0_1(isu__T_284_0_1),
    ._T_284_0_2(isu__T_284_0_2),
    ._T_284_0_3(isu__T_284_0_3),
    ._T_284_0_4(isu__T_284_0_4),
    ._T_284_0_5(isu__T_284_0_5),
    ._T_284_0_6(isu__T_284_0_6),
    ._T_284_0_7(isu__T_284_0_7),
    ._T_284_0_8(isu__T_284_0_8),
    ._T_284_0_9(isu__T_284_0_9),
    ._T_284_0_10(isu__T_284_0_10),
    ._T_284_0_11(isu__T_284_0_11),
    ._T_284_0_12(isu__T_284_0_12),
    ._T_284_0_13(isu__T_284_0_13),
    ._T_284_0_14(isu__T_284_0_14),
    ._T_284_0_15(isu__T_284_0_15),
    ._T_284_0_16(isu__T_284_0_16),
    ._T_284_0_17(isu__T_284_0_17),
    ._T_284_0_18(isu__T_284_0_18),
    ._T_284_0_19(isu__T_284_0_19),
    ._T_284_0_20(isu__T_284_0_20),
    ._T_284_0_21(isu__T_284_0_21),
    ._T_284_0_22(isu__T_284_0_22),
    ._T_284_0_23(isu__T_284_0_23),
    ._T_284_0_24(isu__T_284_0_24),
    ._T_284_0_25(isu__T_284_0_25),
    ._T_284_0_26(isu__T_284_0_26),
    ._T_284_0_27(isu__T_284_0_27),
    ._T_284_0_28(isu__T_284_0_28),
    ._T_284_0_29(isu__T_284_0_29),
    ._T_284_0_30(isu__T_284_0_30),
    ._T_284_0_31(isu__T_284_0_31),
    ._T_186_0(isu__T_186_0),
    .DISPLAY_ENABLE(isu_DISPLAY_ENABLE),
    ._T_187_0(isu__T_187_0)
  );
  EXU exu ( // @[Backend.scala 677:20]
    .clock(exu_clock),
    .reset(exu_reset),
    .io__in_ready(exu_io__in_ready),
    .io__in_valid(exu_io__in_valid),
    .io__in_bits_cf_instr(exu_io__in_bits_cf_instr),
    .io__in_bits_cf_pc(exu_io__in_bits_cf_pc),
    .io__in_bits_cf_pnpc(exu_io__in_bits_cf_pnpc),
    .io__in_bits_cf_exceptionVec_1(exu_io__in_bits_cf_exceptionVec_1),
    .io__in_bits_cf_exceptionVec_2(exu_io__in_bits_cf_exceptionVec_2),
    .io__in_bits_cf_exceptionVec_12(exu_io__in_bits_cf_exceptionVec_12),
    .io__in_bits_cf_intrVec_0(exu_io__in_bits_cf_intrVec_0),
    .io__in_bits_cf_intrVec_1(exu_io__in_bits_cf_intrVec_1),
    .io__in_bits_cf_intrVec_2(exu_io__in_bits_cf_intrVec_2),
    .io__in_bits_cf_intrVec_3(exu_io__in_bits_cf_intrVec_3),
    .io__in_bits_cf_intrVec_4(exu_io__in_bits_cf_intrVec_4),
    .io__in_bits_cf_intrVec_5(exu_io__in_bits_cf_intrVec_5),
    .io__in_bits_cf_intrVec_6(exu_io__in_bits_cf_intrVec_6),
    .io__in_bits_cf_intrVec_7(exu_io__in_bits_cf_intrVec_7),
    .io__in_bits_cf_intrVec_8(exu_io__in_bits_cf_intrVec_8),
    .io__in_bits_cf_intrVec_9(exu_io__in_bits_cf_intrVec_9),
    .io__in_bits_cf_intrVec_10(exu_io__in_bits_cf_intrVec_10),
    .io__in_bits_cf_intrVec_11(exu_io__in_bits_cf_intrVec_11),
    .io__in_bits_cf_brIdx(exu_io__in_bits_cf_brIdx),
    .io__in_bits_cf_crossPageIPFFix(exu_io__in_bits_cf_crossPageIPFFix),
    .io__in_bits_ctrl_fuType(exu_io__in_bits_ctrl_fuType),
    .io__in_bits_ctrl_fuOpType(exu_io__in_bits_ctrl_fuOpType),
    .io__in_bits_ctrl_rfWen(exu_io__in_bits_ctrl_rfWen),
    .io__in_bits_ctrl_rfDest(exu_io__in_bits_ctrl_rfDest),
    .io__in_bits_ctrl_isNutCoreTrap(exu_io__in_bits_ctrl_isNutCoreTrap),
    .io__in_bits_data_src1(exu_io__in_bits_data_src1),
    .io__in_bits_data_src2(exu_io__in_bits_data_src2),
    .io__in_bits_data_imm(exu_io__in_bits_data_imm),
    .io__in_bits_data_srf_0(exu_io__in_bits_data_srf_0),
    .io__in_bits_data_srf_1(exu_io__in_bits_data_srf_1),
    .io__in_bits_data_srf_2(exu_io__in_bits_data_srf_2),
    .io__in_bits_data_srf_3(exu_io__in_bits_data_srf_3),
    .io__out_ready(exu_io__out_ready),
    .io__out_valid(exu_io__out_valid),
    .io__out_bits_decode_cf_instr(exu_io__out_bits_decode_cf_instr),
    .io__out_bits_decode_cf_pc(exu_io__out_bits_decode_cf_pc),
    .io__out_bits_decode_cf_redirect_target(exu_io__out_bits_decode_cf_redirect_target),
    .io__out_bits_decode_cf_redirect_valid(exu_io__out_bits_decode_cf_redirect_valid),
    .io__out_bits_decode_ctrl_fuType(exu_io__out_bits_decode_ctrl_fuType),
    .io__out_bits_decode_ctrl_rfWen(exu_io__out_bits_decode_ctrl_rfWen),
    .io__out_bits_decode_ctrl_rfDest(exu_io__out_bits_decode_ctrl_rfDest),
    .io__out_bits_decode_ctrl_srfWen(exu_io__out_bits_decode_ctrl_srfWen),
    .io__out_bits_decode_ctrl_srfDest(exu_io__out_bits_decode_ctrl_srfDest),
    .io__out_bits_isMMIO(exu_io__out_bits_isMMIO),
    .io__out_bits_intrNO(exu_io__out_bits_intrNO),
    .io__out_bits_commits_0(exu_io__out_bits_commits_0),
    .io__out_bits_commits_1(exu_io__out_bits_commits_1),
    .io__out_bits_commits_2(exu_io__out_bits_commits_2),
    .io__out_bits_commits_3(exu_io__out_bits_commits_3),
    .io__out_bits_commits_5(exu_io__out_bits_commits_5),
    .io__flush(exu_io__flush),
    .io__dmem_req_ready(exu_io__dmem_req_ready),
    .io__dmem_req_valid(exu_io__dmem_req_valid),
    .io__dmem_req_bits_addr(exu_io__dmem_req_bits_addr),
    .io__dmem_req_bits_size(exu_io__dmem_req_bits_size),
    .io__dmem_req_bits_cmd(exu_io__dmem_req_bits_cmd),
    .io__dmem_req_bits_wmask(exu_io__dmem_req_bits_wmask),
    .io__dmem_req_bits_wdata(exu_io__dmem_req_bits_wdata),
    .io__dmem_resp_valid(exu_io__dmem_resp_valid),
    .io__dmem_resp_bits_rdata(exu_io__dmem_resp_bits_rdata),
    .io__forward_valid(exu_io__forward_valid),
    .io__forward_wb_rfWen(exu_io__forward_wb_rfWen),
    .io__forward_wb_rfDest(exu_io__forward_wb_rfDest),
    .io__forward_wb_rfData(exu_io__forward_wb_rfData),
    .io__forward_wb_srfDest(exu_io__forward_wb_srfDest),
    .io__forward_wb_srfData(exu_io__forward_wb_srfData),
    .io__forward_fuType(exu_io__forward_fuType),
    .io__memMMU_imem_priviledgeMode(exu_io__memMMU_imem_priviledgeMode),
    .io__memMMU_dmem_priviledgeMode(exu_io__memMMU_dmem_priviledgeMode),
    .io__memMMU_dmem_status_sum(exu_io__memMMU_dmem_status_sum),
    .io__memMMU_dmem_status_mxr(exu_io__memMMU_dmem_status_mxr),
    .io__memMMU_dmem_loadPF(exu_io__memMMU_dmem_loadPF),
    .io__memMMU_dmem_storePF(exu_io__memMMU_dmem_storePF),
    .io__memMMU_dmem_addr(exu_io__memMMU_dmem_addr),
    ._T_4181(exu__T_4181),
    ._T_4184(exu__T_4184),
    ._T_183(exu__T_183),
    ._T_38_0(exu__T_38_0),
    .flushICache(exu_flushICache),
    ._T_4185(exu__T_4185),
    .satp(exu_satp),
    ._T_243_valid(exu__T_243_valid),
    ._T_243_pc(exu__T_243_pc),
    ._T_243_isMissPredict(exu__T_243_isMissPredict),
    ._T_243_actualTarget(exu__T_243_actualTarget),
    ._T_243_actualTaken(exu__T_243_actualTaken),
    ._T_243_fuOpType(exu__T_243_fuOpType),
    ._T_243_btbType(exu__T_243_btbType),
    ._T_243_isRVC(exu__T_243_isRVC),
    ._T_4178(exu__T_4178),
    .io_in_valid(exu_io_in_valid),
    .mmio(exu_mmio),
    ._T_186(exu__T_186),
    .io_extra_mtip(exu_io_extra_mtip),
    .amoReq(exu_amoReq),
    .DISPLAY_ENABLE(exu_DISPLAY_ENABLE),
    .io_extra_meip_0(exu_io_extra_meip_0),
    ._T_187(exu__T_187),
    .vmEnable(exu_vmEnable),
    .intrVec(exu_intrVec),
    ._T_37_1(exu__T_37_1),
    .io_extra_msip(exu_io_extra_msip),
    ._T_65_0(exu__T_65_0),
    ._T_4183(exu__T_4183),
    ._T_4182(exu__T_4182),
    .flushTLB(exu_flushTLB),
    ._T_66_0(exu__T_66_0),
    ._T_4179(exu__T_4179),
    .falseWire_1(exu_falseWire_1)
  );
  WBU wbu ( // @[Backend.scala 678:20]
    .clock(wbu_clock),
    .reset(wbu_reset),
    .io__in_valid(wbu_io__in_valid),
    .io__in_bits_decode_cf_instr(wbu_io__in_bits_decode_cf_instr),
    .io__in_bits_decode_cf_pc(wbu_io__in_bits_decode_cf_pc),
    .io__in_bits_decode_cf_redirect_target(wbu_io__in_bits_decode_cf_redirect_target),
    .io__in_bits_decode_cf_redirect_valid(wbu_io__in_bits_decode_cf_redirect_valid),
    .io__in_bits_decode_ctrl_fuType(wbu_io__in_bits_decode_ctrl_fuType),
    .io__in_bits_decode_ctrl_rfWen(wbu_io__in_bits_decode_ctrl_rfWen),
    .io__in_bits_decode_ctrl_rfDest(wbu_io__in_bits_decode_ctrl_rfDest),
    .io__in_bits_decode_ctrl_srfWen(wbu_io__in_bits_decode_ctrl_srfWen),
    .io__in_bits_decode_ctrl_srfDest(wbu_io__in_bits_decode_ctrl_srfDest),
    .io__in_bits_isMMIO(wbu_io__in_bits_isMMIO),
    .io__in_bits_intrNO(wbu_io__in_bits_intrNO),
    .io__in_bits_commits_0(wbu_io__in_bits_commits_0),
    .io__in_bits_commits_1(wbu_io__in_bits_commits_1),
    .io__in_bits_commits_2(wbu_io__in_bits_commits_2),
    .io__in_bits_commits_3(wbu_io__in_bits_commits_3),
    .io__in_bits_commits_5(wbu_io__in_bits_commits_5),
    .io__wb_rfWen(wbu_io__wb_rfWen),
    .io__wb_rfDest(wbu_io__wb_rfDest),
    .io__wb_rfData(wbu_io__wb_rfData),
    .io__wb_srfWen(wbu_io__wb_srfWen),
    .io__wb_srfDest(wbu_io__wb_srfDest),
    .io__wb_srfData(wbu_io__wb_srfData),
    .io__redirect_target(wbu_io__redirect_target),
    .io__redirect_valid(wbu_io__redirect_valid),
    .falseWire_0(wbu_falseWire_0),
    .falseWire_1(wbu_falseWire_1),
    .io_in_valid(wbu_io_in_valid),
    ._T_36_0(wbu__T_36_0),
    ._T_32_0(wbu__T_32_0),
    .DISPLAY_ENABLE(wbu_DISPLAY_ENABLE),
    ._T_31_0(wbu__T_31_0),
    ._T_37_0(wbu__T_37_0),
    ._T_26_0(wbu__T_26_0),
    ._T_33_0(wbu__T_33_0),
    .falseWire_2(wbu_falseWire_2)
  );
  assign io_in_0_ready = isu_io_in_0_ready; // @[Backend.scala 683:13]
  assign io_dmem_req_valid = exu_io__dmem_req_valid; // @[Backend.scala 695:11]
  assign io_dmem_req_bits_addr = exu_io__dmem_req_bits_addr; // @[Backend.scala 695:11]
  assign io_dmem_req_bits_size = exu_io__dmem_req_bits_size; // @[Backend.scala 695:11]
  assign io_dmem_req_bits_cmd = exu_io__dmem_req_bits_cmd; // @[Backend.scala 695:11]
  assign io_dmem_req_bits_wmask = exu_io__dmem_req_bits_wmask; // @[Backend.scala 695:11]
  assign io_dmem_req_bits_wdata = exu_io__dmem_req_bits_wdata; // @[Backend.scala 695:11]
  assign io_memMMU_imem_priviledgeMode = exu_io__memMMU_imem_priviledgeMode; // @[Backend.scala 693:18]
  assign io_memMMU_dmem_priviledgeMode = exu_io__memMMU_dmem_priviledgeMode; // @[Backend.scala 694:18]
  assign io_memMMU_dmem_status_sum = exu_io__memMMU_dmem_status_sum; // @[Backend.scala 694:18]
  assign io_memMMU_dmem_status_mxr = exu_io__memMMU_dmem_status_mxr; // @[Backend.scala 694:18]
  assign io_redirect_target = wbu_io__redirect_target; // @[Backend.scala 689:15]
  assign io_redirect_valid = wbu_io__redirect_valid; // @[Backend.scala 689:15]
  assign _T_4181 = exu__T_4181;
  assign _T_4184 = exu__T_4184;
  assign flushICache = exu_flushICache;
  assign _T_4185 = exu__T_4185;
  assign falseWire = wbu_falseWire_0;
  assign satp = exu_satp;
  assign _T_243_valid = exu__T_243_valid;
  assign _T_243_pc = exu__T_243_pc;
  assign _T_243_isMissPredict = exu__T_243_isMissPredict;
  assign _T_243_actualTarget = exu__T_243_actualTarget;
  assign _T_243_actualTaken = exu__T_243_actualTaken;
  assign _T_243_fuOpType = exu__T_243_fuOpType;
  assign _T_243_btbType = exu__T_243_btbType;
  assign _T_243_isRVC = exu__T_243_isRVC;
  assign falseWire_0 = wbu_falseWire_1;
  assign _T_4178 = exu__T_4178;
  assign _T_284_0 = isu__T_284_0_0;
  assign _T_284_1 = isu__T_284_0_1;
  assign _T_284_2 = isu__T_284_0_2;
  assign _T_284_3 = isu__T_284_0_3;
  assign _T_284_4 = isu__T_284_0_4;
  assign _T_284_5 = isu__T_284_0_5;
  assign _T_284_6 = isu__T_284_0_6;
  assign _T_284_7 = isu__T_284_0_7;
  assign _T_284_8 = isu__T_284_0_8;
  assign _T_284_9 = isu__T_284_0_9;
  assign _T_284_10 = isu__T_284_0_10;
  assign _T_284_11 = isu__T_284_0_11;
  assign _T_284_12 = isu__T_284_0_12;
  assign _T_284_13 = isu__T_284_0_13;
  assign _T_284_14 = isu__T_284_0_14;
  assign _T_284_15 = isu__T_284_0_15;
  assign _T_284_16 = isu__T_284_0_16;
  assign _T_284_17 = isu__T_284_0_17;
  assign _T_284_18 = isu__T_284_0_18;
  assign _T_284_19 = isu__T_284_0_19;
  assign _T_284_20 = isu__T_284_0_20;
  assign _T_284_21 = isu__T_284_0_21;
  assign _T_284_22 = isu__T_284_0_22;
  assign _T_284_23 = isu__T_284_0_23;
  assign _T_284_24 = isu__T_284_0_24;
  assign _T_284_25 = isu__T_284_0_25;
  assign _T_284_26 = isu__T_284_0_26;
  assign _T_284_27 = isu__T_284_0_27;
  assign _T_284_28 = isu__T_284_0_28;
  assign _T_284_29 = isu__T_284_0_29;
  assign _T_284_30 = isu__T_284_0_30;
  assign _T_284_31 = isu__T_284_0_31;
  assign _T_36 = wbu__T_36_0;
  assign amoReq = exu_amoReq;
  assign _T_32 = wbu__T_32_0;
  assign _T_31 = wbu__T_31_0;
  assign _T_37 = wbu__T_37_0;
  assign _T_26 = wbu__T_26_0;
  assign intrVec = exu_intrVec;
  assign _T_4183 = exu__T_4183;
  assign _T_4182 = exu__T_4182;
  assign flushTLB = exu_flushTLB;
  assign _T_33 = wbu__T_33_0;
  assign _T_4179 = exu__T_4179;
  assign isu_clock = clock;
  assign isu_reset = reset;
  assign isu_io_in_0_valid = io_in_0_valid; // @[Backend.scala 683:13]
  assign isu_io_in_0_bits_cf_instr = io_in_0_bits_cf_instr; // @[Backend.scala 683:13]
  assign isu_io_in_0_bits_cf_pc = io_in_0_bits_cf_pc; // @[Backend.scala 683:13]
  assign isu_io_in_0_bits_cf_pnpc = io_in_0_bits_cf_pnpc; // @[Backend.scala 683:13]
  assign isu_io_in_0_bits_cf_exceptionVec_1 = io_in_0_bits_cf_exceptionVec_1; // @[Backend.scala 683:13]
  assign isu_io_in_0_bits_cf_exceptionVec_2 = io_in_0_bits_cf_exceptionVec_2; // @[Backend.scala 683:13]
  assign isu_io_in_0_bits_cf_exceptionVec_12 = io_in_0_bits_cf_exceptionVec_12; // @[Backend.scala 683:13]
  assign isu_io_in_0_bits_cf_intrVec_0 = io_in_0_bits_cf_intrVec_0; // @[Backend.scala 683:13]
  assign isu_io_in_0_bits_cf_intrVec_1 = io_in_0_bits_cf_intrVec_1; // @[Backend.scala 683:13]
  assign isu_io_in_0_bits_cf_intrVec_2 = io_in_0_bits_cf_intrVec_2; // @[Backend.scala 683:13]
  assign isu_io_in_0_bits_cf_intrVec_3 = io_in_0_bits_cf_intrVec_3; // @[Backend.scala 683:13]
  assign isu_io_in_0_bits_cf_intrVec_4 = io_in_0_bits_cf_intrVec_4; // @[Backend.scala 683:13]
  assign isu_io_in_0_bits_cf_intrVec_5 = io_in_0_bits_cf_intrVec_5; // @[Backend.scala 683:13]
  assign isu_io_in_0_bits_cf_intrVec_6 = io_in_0_bits_cf_intrVec_6; // @[Backend.scala 683:13]
  assign isu_io_in_0_bits_cf_intrVec_7 = io_in_0_bits_cf_intrVec_7; // @[Backend.scala 683:13]
  assign isu_io_in_0_bits_cf_intrVec_8 = io_in_0_bits_cf_intrVec_8; // @[Backend.scala 683:13]
  assign isu_io_in_0_bits_cf_intrVec_9 = io_in_0_bits_cf_intrVec_9; // @[Backend.scala 683:13]
  assign isu_io_in_0_bits_cf_intrVec_10 = io_in_0_bits_cf_intrVec_10; // @[Backend.scala 683:13]
  assign isu_io_in_0_bits_cf_intrVec_11 = io_in_0_bits_cf_intrVec_11; // @[Backend.scala 683:13]
  assign isu_io_in_0_bits_cf_brIdx = io_in_0_bits_cf_brIdx; // @[Backend.scala 683:13]
  assign isu_io_in_0_bits_cf_crossPageIPFFix = io_in_0_bits_cf_crossPageIPFFix; // @[Backend.scala 683:13]
  assign isu_io_in_0_bits_ctrl_src1Type = io_in_0_bits_ctrl_src1Type; // @[Backend.scala 683:13]
  assign isu_io_in_0_bits_ctrl_src2Type = io_in_0_bits_ctrl_src2Type; // @[Backend.scala 683:13]
  assign isu_io_in_0_bits_ctrl_fuType = io_in_0_bits_ctrl_fuType; // @[Backend.scala 683:13]
  assign isu_io_in_0_bits_ctrl_fuOpType = io_in_0_bits_ctrl_fuOpType; // @[Backend.scala 683:13]
  assign isu_io_in_0_bits_ctrl_rfSrc1 = io_in_0_bits_ctrl_rfSrc1; // @[Backend.scala 683:13]
  assign isu_io_in_0_bits_ctrl_rfSrc2 = io_in_0_bits_ctrl_rfSrc2; // @[Backend.scala 683:13]
  assign isu_io_in_0_bits_ctrl_rfWen = io_in_0_bits_ctrl_rfWen; // @[Backend.scala 683:13]
  assign isu_io_in_0_bits_ctrl_rfDest = io_in_0_bits_ctrl_rfDest; // @[Backend.scala 683:13]
  assign isu_io_in_0_bits_ctrl_isNutCoreTrap = io_in_0_bits_ctrl_isNutCoreTrap; // @[Backend.scala 683:13]
  assign isu_io_in_0_bits_data_imm = io_in_0_bits_data_imm; // @[Backend.scala 683:13]
  assign isu_io_out_ready = exu_io__in_ready; // @[Pipeline.scala 29:16]
  assign isu_io_wb_rfWen = wbu_io__wb_rfWen; // @[Backend.scala 687:13]
  assign isu_io_wb_rfDest = wbu_io__wb_rfDest; // @[Backend.scala 687:13]
  assign isu_io_wb_rfData = wbu_io__wb_rfData; // @[Backend.scala 687:13]
  assign isu_io_wb_srfWen = wbu_io__wb_srfWen; // @[Backend.scala 687:13]
  assign isu_io_wb_srfDest = wbu_io__wb_srfDest; // @[Backend.scala 687:13]
  assign isu_io_wb_srfData = wbu_io__wb_srfData; // @[Backend.scala 687:13]
  assign isu_io_forward_valid = exu_io__forward_valid; // @[Backend.scala 691:18]
  assign isu_io_forward_wb_rfWen = exu_io__forward_wb_rfWen; // @[Backend.scala 691:18]
  assign isu_io_forward_wb_rfDest = exu_io__forward_wb_rfDest; // @[Backend.scala 691:18]
  assign isu_io_forward_wb_rfData = exu_io__forward_wb_rfData; // @[Backend.scala 691:18]
  assign isu_io_forward_wb_srfDest = exu_io__forward_wb_srfDest; // @[Backend.scala 691:18]
  assign isu_io_forward_wb_srfData = exu_io__forward_wb_srfData; // @[Backend.scala 691:18]
  assign isu_io_forward_fuType = exu_io__forward_fuType; // @[Backend.scala 691:18]
  assign isu_io_flush = io_flush[0]; // @[Backend.scala 685:16]
  assign isu_DISPLAY_ENABLE = _T_13;
  assign exu_clock = clock;
  assign exu_reset = reset;
  assign exu_io__in_valid = _T_2; // @[Pipeline.scala 31:17]
  assign exu_io__in_bits_cf_instr = _T_5_cf_instr; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_pc = _T_5_cf_pc; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_pnpc = _T_5_cf_pnpc; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_exceptionVec_1 = _T_5_cf_exceptionVec_1; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_exceptionVec_2 = _T_5_cf_exceptionVec_2; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_exceptionVec_12 = _T_5_cf_exceptionVec_12; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_0 = _T_5_cf_intrVec_0; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_1 = _T_5_cf_intrVec_1; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_2 = _T_5_cf_intrVec_2; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_3 = _T_5_cf_intrVec_3; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_4 = _T_5_cf_intrVec_4; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_5 = _T_5_cf_intrVec_5; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_6 = _T_5_cf_intrVec_6; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_7 = _T_5_cf_intrVec_7; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_8 = _T_5_cf_intrVec_8; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_9 = _T_5_cf_intrVec_9; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_10 = _T_5_cf_intrVec_10; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_11 = _T_5_cf_intrVec_11; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_brIdx = _T_5_cf_brIdx; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_crossPageIPFFix = _T_5_cf_crossPageIPFFix; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_fuType = _T_5_ctrl_fuType; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_fuOpType = _T_5_ctrl_fuOpType; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_rfWen = _T_5_ctrl_rfWen; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_rfDest = _T_5_ctrl_rfDest; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_isNutCoreTrap = _T_5_ctrl_isNutCoreTrap; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_data_src1 = _T_5_data_src1; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_data_src2 = _T_5_data_src2; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_data_imm = _T_5_data_imm; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_data_srf_0 = _T_5_data_srf_0; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_data_srf_1 = _T_5_data_srf_1; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_data_srf_2 = _T_5_data_srf_2; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_data_srf_3 = _T_5_data_srf_3; // @[Pipeline.scala 30:16]
  assign exu_io__out_ready = 1'h1; // @[Pipeline.scala 29:16]
  assign exu_io__flush = io_flush[1]; // @[Backend.scala 686:16]
  assign exu_io__dmem_req_ready = io_dmem_req_ready; // @[Backend.scala 695:11]
  assign exu_io__dmem_resp_valid = io_dmem_resp_valid; // @[Backend.scala 695:11]
  assign exu_io__dmem_resp_bits_rdata = io_dmem_resp_bits_rdata; // @[Backend.scala 695:11]
  assign exu_io__memMMU_dmem_loadPF = io_memMMU_dmem_loadPF; // @[Backend.scala 694:18]
  assign exu_io__memMMU_dmem_storePF = io_memMMU_dmem_storePF; // @[Backend.scala 694:18]
  assign exu_io__memMMU_dmem_addr = io_memMMU_dmem_addr; // @[Backend.scala 694:18]
  assign exu__T_183 = isu__T_183_0;
  assign exu__T_38_0 = _T_38;
  assign exu_io_in_valid = wbu_io_in_valid;
  assign exu_mmio = mmio;
  assign exu__T_186 = isu__T_186_0;
  assign exu_io_extra_mtip = io_extra_mtip;
  assign exu_DISPLAY_ENABLE = _T_13;
  assign exu_io_extra_meip_0 = io_extra_meip_0;
  assign exu__T_187 = isu__T_187_0;
  assign exu_vmEnable = vmEnable;
  assign exu__T_37_1 = _T_37_0;
  assign exu_io_extra_msip = io_extra_msip;
  assign exu__T_65_0 = _T_65;
  assign exu__T_66_0 = _T_66;
  assign exu_falseWire_1 = wbu_falseWire_2;
  assign wbu_clock = clock;
  assign wbu_reset = reset;
  assign wbu_io__in_valid = _T_7; // @[Pipeline.scala 31:17]
  assign wbu_io__in_bits_decode_cf_instr = _T_10_decode_cf_instr; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_cf_pc = _T_10_decode_cf_pc; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_cf_redirect_target = _T_10_decode_cf_redirect_target; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_cf_redirect_valid = _T_10_decode_cf_redirect_valid; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_ctrl_fuType = _T_10_decode_ctrl_fuType; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_ctrl_rfWen = _T_10_decode_ctrl_rfWen; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_ctrl_rfDest = _T_10_decode_ctrl_rfDest; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_ctrl_srfWen = _T_10_decode_ctrl_srfWen; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_ctrl_srfDest = _T_10_decode_ctrl_srfDest; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_isMMIO = _T_10_isMMIO; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_intrNO = _T_10_intrNO; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_0 = _T_10_commits_0; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_1 = _T_10_commits_1; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_2 = _T_10_commits_2; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_3 = _T_10_commits_3; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_5 = _T_10_commits_5; // @[Pipeline.scala 30:16]
  assign wbu_DISPLAY_ENABLE = _T_13;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_2 = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  _T_5_cf_instr = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  _T_5_cf_pc = _RAND_2[38:0];
  _RAND_3 = {2{`RANDOM}};
  _T_5_cf_pnpc = _RAND_3[38:0];
  _RAND_4 = {1{`RANDOM}};
  _T_5_cf_exceptionVec_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _T_5_cf_exceptionVec_2 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _T_5_cf_exceptionVec_12 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_5_cf_intrVec_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _T_5_cf_intrVec_1 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _T_5_cf_intrVec_2 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _T_5_cf_intrVec_3 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _T_5_cf_intrVec_4 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _T_5_cf_intrVec_5 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _T_5_cf_intrVec_6 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  _T_5_cf_intrVec_7 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  _T_5_cf_intrVec_8 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  _T_5_cf_intrVec_9 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  _T_5_cf_intrVec_10 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  _T_5_cf_intrVec_11 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  _T_5_cf_brIdx = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  _T_5_cf_crossPageIPFFix = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  _T_5_ctrl_fuType = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  _T_5_ctrl_fuOpType = _RAND_22[6:0];
  _RAND_23 = {1{`RANDOM}};
  _T_5_ctrl_rfWen = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  _T_5_ctrl_rfDest = _RAND_24[4:0];
  _RAND_25 = {1{`RANDOM}};
  _T_5_ctrl_isNutCoreTrap = _RAND_25[0:0];
  _RAND_26 = {2{`RANDOM}};
  _T_5_data_src1 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  _T_5_data_src2 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  _T_5_data_imm = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  _T_5_data_srf_0 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  _T_5_data_srf_1 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  _T_5_data_srf_2 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  _T_5_data_srf_3 = _RAND_32[63:0];
  _RAND_33 = {1{`RANDOM}};
  _T_7 = _RAND_33[0:0];
  _RAND_34 = {2{`RANDOM}};
  _T_10_decode_cf_instr = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  _T_10_decode_cf_pc = _RAND_35[38:0];
  _RAND_36 = {2{`RANDOM}};
  _T_10_decode_cf_redirect_target = _RAND_36[38:0];
  _RAND_37 = {1{`RANDOM}};
  _T_10_decode_cf_redirect_valid = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  _T_10_decode_ctrl_fuType = _RAND_38[2:0];
  _RAND_39 = {1{`RANDOM}};
  _T_10_decode_ctrl_rfWen = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  _T_10_decode_ctrl_rfDest = _RAND_40[4:0];
  _RAND_41 = {1{`RANDOM}};
  _T_10_decode_ctrl_srfWen = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  _T_10_decode_ctrl_srfDest = _RAND_42[2:0];
  _RAND_43 = {1{`RANDOM}};
  _T_10_isMMIO = _RAND_43[0:0];
  _RAND_44 = {2{`RANDOM}};
  _T_10_intrNO = _RAND_44[63:0];
  _RAND_45 = {2{`RANDOM}};
  _T_10_commits_0 = _RAND_45[63:0];
  _RAND_46 = {2{`RANDOM}};
  _T_10_commits_1 = _RAND_46[63:0];
  _RAND_47 = {2{`RANDOM}};
  _T_10_commits_2 = _RAND_47[63:0];
  _RAND_48 = {2{`RANDOM}};
  _T_10_commits_3 = _RAND_48[63:0];
  _RAND_49 = {2{`RANDOM}};
  _T_10_commits_5 = _RAND_49[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_2 <= 1'h0;
    end else if (io_flush[0]) begin
      _T_2 <= 1'h0;
    end else begin
      _T_2 <= _GEN_1;
    end
    if (_T_3) begin
      _T_5_cf_instr <= isu_io_out_bits_cf_instr;
    end
    if (_T_3) begin
      _T_5_cf_pc <= isu_io_out_bits_cf_pc;
    end
    if (_T_3) begin
      _T_5_cf_pnpc <= isu_io_out_bits_cf_pnpc;
    end
    if (_T_3) begin
      _T_5_cf_exceptionVec_1 <= isu_io_out_bits_cf_exceptionVec_1;
    end
    if (_T_3) begin
      _T_5_cf_exceptionVec_2 <= isu_io_out_bits_cf_exceptionVec_2;
    end
    if (_T_3) begin
      _T_5_cf_exceptionVec_12 <= isu_io_out_bits_cf_exceptionVec_12;
    end
    if (_T_3) begin
      _T_5_cf_intrVec_0 <= isu_io_out_bits_cf_intrVec_0;
    end
    if (_T_3) begin
      _T_5_cf_intrVec_1 <= isu_io_out_bits_cf_intrVec_1;
    end
    if (_T_3) begin
      _T_5_cf_intrVec_2 <= isu_io_out_bits_cf_intrVec_2;
    end
    if (_T_3) begin
      _T_5_cf_intrVec_3 <= isu_io_out_bits_cf_intrVec_3;
    end
    if (_T_3) begin
      _T_5_cf_intrVec_4 <= isu_io_out_bits_cf_intrVec_4;
    end
    if (_T_3) begin
      _T_5_cf_intrVec_5 <= isu_io_out_bits_cf_intrVec_5;
    end
    if (_T_3) begin
      _T_5_cf_intrVec_6 <= isu_io_out_bits_cf_intrVec_6;
    end
    if (_T_3) begin
      _T_5_cf_intrVec_7 <= isu_io_out_bits_cf_intrVec_7;
    end
    if (_T_3) begin
      _T_5_cf_intrVec_8 <= isu_io_out_bits_cf_intrVec_8;
    end
    if (_T_3) begin
      _T_5_cf_intrVec_9 <= isu_io_out_bits_cf_intrVec_9;
    end
    if (_T_3) begin
      _T_5_cf_intrVec_10 <= isu_io_out_bits_cf_intrVec_10;
    end
    if (_T_3) begin
      _T_5_cf_intrVec_11 <= isu_io_out_bits_cf_intrVec_11;
    end
    if (_T_3) begin
      _T_5_cf_brIdx <= isu_io_out_bits_cf_brIdx;
    end
    if (_T_3) begin
      _T_5_cf_crossPageIPFFix <= isu_io_out_bits_cf_crossPageIPFFix;
    end
    if (_T_3) begin
      _T_5_ctrl_fuType <= isu_io_out_bits_ctrl_fuType;
    end
    if (_T_3) begin
      _T_5_ctrl_fuOpType <= isu_io_out_bits_ctrl_fuOpType;
    end
    if (_T_3) begin
      _T_5_ctrl_rfWen <= isu_io_out_bits_ctrl_rfWen;
    end
    if (_T_3) begin
      _T_5_ctrl_rfDest <= isu_io_out_bits_ctrl_rfDest;
    end
    if (_T_3) begin
      _T_5_ctrl_isNutCoreTrap <= isu_io_out_bits_ctrl_isNutCoreTrap;
    end
    if (_T_3) begin
      _T_5_data_src1 <= isu_io_out_bits_data_src1;
    end
    if (_T_3) begin
      _T_5_data_src2 <= isu_io_out_bits_data_src2;
    end
    if (_T_3) begin
      _T_5_data_imm <= isu_io_out_bits_data_imm;
    end
    if (_T_3) begin
      _T_5_data_srf_0 <= isu_io_out_bits_data_srf_0;
    end
    if (_T_3) begin
      _T_5_data_srf_1 <= isu_io_out_bits_data_srf_1;
    end
    if (_T_3) begin
      _T_5_data_srf_2 <= isu_io_out_bits_data_srf_2;
    end
    if (_T_3) begin
      _T_5_data_srf_3 <= isu_io_out_bits_data_srf_3;
    end
    if (reset) begin
      _T_7 <= 1'h0;
    end else if (io_flush[1]) begin
      _T_7 <= 1'h0;
    end else begin
      _T_7 <= _T_8;
    end
    if (_T_8) begin
      _T_10_decode_cf_instr <= exu_io__out_bits_decode_cf_instr;
    end
    if (_T_8) begin
      _T_10_decode_cf_pc <= exu_io__out_bits_decode_cf_pc;
    end
    if (_T_8) begin
      _T_10_decode_cf_redirect_target <= exu_io__out_bits_decode_cf_redirect_target;
    end
    if (_T_8) begin
      _T_10_decode_cf_redirect_valid <= exu_io__out_bits_decode_cf_redirect_valid;
    end
    if (_T_8) begin
      _T_10_decode_ctrl_fuType <= exu_io__out_bits_decode_ctrl_fuType;
    end
    if (_T_8) begin
      _T_10_decode_ctrl_rfWen <= exu_io__out_bits_decode_ctrl_rfWen;
    end
    if (_T_8) begin
      _T_10_decode_ctrl_rfDest <= exu_io__out_bits_decode_ctrl_rfDest;
    end
    if (_T_8) begin
      _T_10_decode_ctrl_srfWen <= exu_io__out_bits_decode_ctrl_srfWen;
    end
    if (_T_8) begin
      _T_10_decode_ctrl_srfDest <= exu_io__out_bits_decode_ctrl_srfDest;
    end
    if (_T_8) begin
      _T_10_isMMIO <= exu_io__out_bits_isMMIO;
    end
    if (_T_8) begin
      _T_10_intrNO <= exu_io__out_bits_intrNO;
    end
    if (_T_8) begin
      _T_10_commits_0 <= exu_io__out_bits_commits_0;
    end
    if (_T_8) begin
      _T_10_commits_1 <= exu_io__out_bits_commits_1;
    end
    if (_T_8) begin
      _T_10_commits_2 <= exu_io__out_bits_commits_2;
    end
    if (_T_8) begin
      _T_10_commits_3 <= exu_io__out_bits_commits_3;
    end
    if (_T_8) begin
      _T_10_commits_5 <= exu_io__out_bits_commits_5;
    end
  end
endmodule
module LockingArbiter(
  input         clock,
  input         reset,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input  [3:0]  io_in_0_bits_cmd,
  input  [7:0]  io_in_0_bits_wmask,
  input  [63:0] io_in_0_bits_wdata,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input  [2:0]  io_in_1_bits_size,
  input  [3:0]  io_in_1_bits_cmd,
  input  [7:0]  io_in_1_bits_wmask,
  input  [63:0] io_in_1_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [2:0]  io_out_bits_size,
  output [3:0]  io_out_bits_cmd,
  output [7:0]  io_out_bits_wmask,
  output [63:0] io_out_bits_wdata,
  output        io_chosen
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] value; // @[Counter.scala 29:33]
  reg  _T; // @[Arbiter.scala 46:22]
  wire  _T_1 = value != 3'h0; // @[Arbiter.scala 47:34]
  wire  _T_4 = io_out_bits_cmd[0] & io_out_bits_cmd[1]; // @[Crossbar.scala 100:62]
  wire  _T_5 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_6 = _T_5 & _T_4; // @[Arbiter.scala 50:25]
  wire [2:0] _T_9 = value + 3'h1; // @[Counter.scala 39:22]
  wire  choice = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbiter.scala 88:27]
  wire  _T_10 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  wire  _T_11 = ~_T; // @[Arbiter.scala 57:39]
  wire  _T_12 = _T_1 ? _T_11 : 1'h1; // @[Arbiter.scala 57:22]
  wire  _T_15 = _T_1 ? _T : _T_10; // @[Arbiter.scala 57:22]
  assign io_in_0_ready = _T_12 & io_out_ready; // @[Arbiter.scala 57:16]
  assign io_in_1_ready = _T_15 & io_out_ready; // @[Arbiter.scala 57:16]
  assign io_out_valid = io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 41:16]
  assign io_out_bits_addr = io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr; // @[Arbiter.scala 42:15]
  assign io_out_bits_size = io_chosen ? io_in_1_bits_size : 3'h3; // @[Arbiter.scala 42:15]
  assign io_out_bits_cmd = io_chosen ? io_in_1_bits_cmd : io_in_0_bits_cmd; // @[Arbiter.scala 42:15]
  assign io_out_bits_wmask = io_chosen ? io_in_1_bits_wmask : io_in_0_bits_wmask; // @[Arbiter.scala 42:15]
  assign io_out_bits_wdata = io_chosen ? io_in_1_bits_wdata : io_in_0_bits_wdata; // @[Arbiter.scala 42:15]
  assign io_chosen = _T_1 ? _T : choice; // @[Arbiter.scala 40:13 Arbiter.scala 55:31]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  _T = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 3'h0;
    end else if (_T_6) begin
      value <= _T_9;
    end
    if (_T_6) begin
      _T <= io_chosen;
    end
  end
endmodule
module SimpleBusCrossbarNto1(
  input         clock,
  input         reset,
  output        io_in_0_req_ready,
  input         io_in_0_req_valid,
  input  [31:0] io_in_0_req_bits_addr,
  input  [3:0]  io_in_0_req_bits_cmd,
  input  [7:0]  io_in_0_req_bits_wmask,
  input  [63:0] io_in_0_req_bits_wdata,
  output        io_in_0_resp_valid,
  output [3:0]  io_in_0_resp_bits_cmd,
  output [63:0] io_in_0_resp_bits_rdata,
  output        io_in_1_req_ready,
  input         io_in_1_req_valid,
  input  [31:0] io_in_1_req_bits_addr,
  input  [2:0]  io_in_1_req_bits_size,
  input  [3:0]  io_in_1_req_bits_cmd,
  input  [7:0]  io_in_1_req_bits_wmask,
  input  [63:0] io_in_1_req_bits_wdata,
  output        io_in_1_resp_valid,
  output [3:0]  io_in_1_resp_bits_cmd,
  output [63:0] io_in_1_resp_bits_rdata,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [2:0]  io_out_req_bits_size,
  output [3:0]  io_out_req_bits_cmd,
  output [7:0]  io_out_req_bits_wmask,
  output [63:0] io_out_req_bits_wdata,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [3:0]  io_out_resp_bits_cmd,
  input  [63:0] io_out_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  inputArb_clock; // @[Crossbar.scala 101:24]
  wire  inputArb_reset; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_0_ready; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_0_valid; // @[Crossbar.scala 101:24]
  wire [31:0] inputArb_io_in_0_bits_addr; // @[Crossbar.scala 101:24]
  wire [3:0] inputArb_io_in_0_bits_cmd; // @[Crossbar.scala 101:24]
  wire [7:0] inputArb_io_in_0_bits_wmask; // @[Crossbar.scala 101:24]
  wire [63:0] inputArb_io_in_0_bits_wdata; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_1_ready; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_1_valid; // @[Crossbar.scala 101:24]
  wire [31:0] inputArb_io_in_1_bits_addr; // @[Crossbar.scala 101:24]
  wire [2:0] inputArb_io_in_1_bits_size; // @[Crossbar.scala 101:24]
  wire [3:0] inputArb_io_in_1_bits_cmd; // @[Crossbar.scala 101:24]
  wire [7:0] inputArb_io_in_1_bits_wmask; // @[Crossbar.scala 101:24]
  wire [63:0] inputArb_io_in_1_bits_wdata; // @[Crossbar.scala 101:24]
  wire  inputArb_io_out_ready; // @[Crossbar.scala 101:24]
  wire  inputArb_io_out_valid; // @[Crossbar.scala 101:24]
  wire [31:0] inputArb_io_out_bits_addr; // @[Crossbar.scala 101:24]
  wire [2:0] inputArb_io_out_bits_size; // @[Crossbar.scala 101:24]
  wire [3:0] inputArb_io_out_bits_cmd; // @[Crossbar.scala 101:24]
  wire [7:0] inputArb_io_out_bits_wmask; // @[Crossbar.scala 101:24]
  wire [63:0] inputArb_io_out_bits_wdata; // @[Crossbar.scala 101:24]
  wire  inputArb_io_chosen; // @[Crossbar.scala 101:24]
  reg [1:0] state; // @[Crossbar.scala 98:22]
  wire  _T_1 = ~inputArb_io_out_bits_cmd[0]; // @[SimpleBus.scala 73:18]
  wire  _T_3 = ~inputArb_io_out_bits_cmd[3]; // @[SimpleBus.scala 73:29]
  wire  _T_4 = _T_1 & _T_3; // @[SimpleBus.scala 73:26]
  wire  _T_5 = ~_T_4; // @[Crossbar.scala 104:29]
  wire  _T_6 = inputArb_io_out_valid & _T_5; // @[Crossbar.scala 104:26]
  wire  _T_9 = _T_6 & _T_1; // @[Crossbar.scala 104:52]
  wire  _T_10 = ~_T_9; // @[Crossbar.scala 104:10]
  wire  _T_12 = _T_10 | reset; // @[Crossbar.scala 104:9]
  wire  _T_13 = ~_T_12; // @[Crossbar.scala 104:9]
  reg  inflightSrc; // @[Crossbar.scala 105:24]
  wire  _T_14 = state == 2'h0; // @[Crossbar.scala 109:47]
  wire  _GEN_34 = ~inflightSrc; // @[Crossbar.scala 115:13]
  wire  _T_18 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_19 = inputArb_io_out_ready & inputArb_io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_25 = inputArb_io_out_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_26 = inputArb_io_out_bits_cmd == 4'h1; // @[SimpleBus.scala 77:29]
  wire  _T_27 = _T_25 | _T_26; // @[Crossbar.scala 124:47]
  wire  _T_28 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_29 = io_out_resp_ready & io_out_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_30 = io_out_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire  _T_31 = _T_29 & _T_30; // @[Crossbar.scala 127:48]
  wire  _T_32 = 2'h2 == state; // @[Conditional.scala 37:30]
  LockingArbiter inputArb ( // @[Crossbar.scala 101:24]
    .clock(inputArb_clock),
    .reset(inputArb_reset),
    .io_in_0_ready(inputArb_io_in_0_ready),
    .io_in_0_valid(inputArb_io_in_0_valid),
    .io_in_0_bits_addr(inputArb_io_in_0_bits_addr),
    .io_in_0_bits_cmd(inputArb_io_in_0_bits_cmd),
    .io_in_0_bits_wmask(inputArb_io_in_0_bits_wmask),
    .io_in_0_bits_wdata(inputArb_io_in_0_bits_wdata),
    .io_in_1_ready(inputArb_io_in_1_ready),
    .io_in_1_valid(inputArb_io_in_1_valid),
    .io_in_1_bits_addr(inputArb_io_in_1_bits_addr),
    .io_in_1_bits_size(inputArb_io_in_1_bits_size),
    .io_in_1_bits_cmd(inputArb_io_in_1_bits_cmd),
    .io_in_1_bits_wmask(inputArb_io_in_1_bits_wmask),
    .io_in_1_bits_wdata(inputArb_io_in_1_bits_wdata),
    .io_out_ready(inputArb_io_out_ready),
    .io_out_valid(inputArb_io_out_valid),
    .io_out_bits_addr(inputArb_io_out_bits_addr),
    .io_out_bits_size(inputArb_io_out_bits_size),
    .io_out_bits_cmd(inputArb_io_out_bits_cmd),
    .io_out_bits_wmask(inputArb_io_out_bits_wmask),
    .io_out_bits_wdata(inputArb_io_out_bits_wdata),
    .io_chosen(inputArb_io_chosen)
  );
  assign io_in_0_req_ready = inputArb_io_in_0_ready; // @[Crossbar.scala 102:68]
  assign io_in_0_resp_valid = _GEN_34 & io_out_resp_valid; // @[Crossbar.scala 113:26 Crossbar.scala 115:13]
  assign io_in_0_resp_bits_cmd = io_out_resp_bits_cmd; // @[Crossbar.scala 112:25]
  assign io_in_0_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 112:25]
  assign io_in_1_req_ready = inputArb_io_in_1_ready; // @[Crossbar.scala 102:68]
  assign io_in_1_resp_valid = inflightSrc & io_out_resp_valid; // @[Crossbar.scala 113:26 Crossbar.scala 115:13]
  assign io_in_1_resp_bits_cmd = io_out_resp_bits_cmd; // @[Crossbar.scala 112:25]
  assign io_in_1_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 112:25]
  assign io_out_req_valid = inputArb_io_out_valid & _T_14; // @[Crossbar.scala 109:20]
  assign io_out_req_bits_addr = inputArb_io_out_bits_addr; // @[Crossbar.scala 107:19]
  assign io_out_req_bits_size = inputArb_io_out_bits_size; // @[Crossbar.scala 107:19]
  assign io_out_req_bits_cmd = inputArb_io_out_bits_cmd; // @[Crossbar.scala 107:19]
  assign io_out_req_bits_wmask = inputArb_io_out_bits_wmask; // @[Crossbar.scala 107:19]
  assign io_out_req_bits_wdata = inputArb_io_out_bits_wdata; // @[Crossbar.scala 107:19]
  assign io_out_resp_ready = 1'h1; // @[Crossbar.scala 116:13]
  assign inputArb_clock = clock;
  assign inputArb_reset = reset;
  assign inputArb_io_in_0_valid = io_in_0_req_valid; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_addr = io_in_0_req_bits_addr; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_cmd = io_in_0_req_bits_cmd; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_wmask = io_in_0_req_bits_wmask; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_wdata = io_in_0_req_bits_wdata; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_valid = io_in_1_req_valid; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_bits_addr = io_in_1_req_bits_addr; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_bits_size = io_in_1_req_bits_size; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_bits_cmd = io_in_1_req_bits_cmd; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_bits_wmask = io_in_1_req_bits_wmask; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_bits_wdata = io_in_1_req_bits_wdata; // @[Crossbar.scala 102:68]
  assign inputArb_io_out_ready = io_out_req_ready & _T_14; // @[Crossbar.scala 110:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  inflightSrc = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else if (_T_18) begin
      if (_T_19) begin
        if (_T_4) begin
          state <= 2'h1;
        end else if (_T_27) begin
          state <= 2'h2;
        end
      end
    end else if (_T_28) begin
      if (_T_31) begin
        state <= 2'h0;
      end
    end else if (_T_32) begin
      if (_T_29) begin
        state <= 2'h0;
      end
    end
    if (_T_18) begin
      if (_T_19) begin
        inflightSrc <= inputArb_io_chosen;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Crossbar.scala:104 assert(!(thisReq.valid && !thisReq.bits.isRead() && !thisReq.bits.isWrite()))\n"); // @[Crossbar.scala 104:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_13) begin
          $fatal; // @[Crossbar.scala 104:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module LockingArbiter_1(
  input         clock,
  input         reset,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input  [2:0]  io_in_0_bits_size,
  input  [3:0]  io_in_0_bits_cmd,
  input  [7:0]  io_in_0_bits_wmask,
  input  [63:0] io_in_0_bits_wdata,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input  [3:0]  io_in_1_bits_cmd,
  input  [63:0] io_in_1_bits_wdata,
  output        io_in_2_ready,
  input         io_in_2_valid,
  input  [31:0] io_in_2_bits_addr,
  input  [3:0]  io_in_2_bits_cmd,
  input  [63:0] io_in_2_bits_wdata,
  output        io_in_3_ready,
  input         io_in_3_valid,
  input  [31:0] io_in_3_bits_addr,
  input  [2:0]  io_in_3_bits_size,
  input  [3:0]  io_in_3_bits_cmd,
  input  [7:0]  io_in_3_bits_wmask,
  input  [63:0] io_in_3_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [2:0]  io_out_bits_size,
  output [3:0]  io_out_bits_cmd,
  output [7:0]  io_out_bits_wmask,
  output [63:0] io_out_bits_wdata,
  output [1:0]  io_chosen
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  _GEN_8 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 41:16]
  wire [31:0] _GEN_9 = 2'h1 == io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr; // @[Arbiter.scala 41:16]
  wire [2:0] _GEN_10 = 2'h1 == io_chosen ? 3'h3 : io_in_0_bits_size; // @[Arbiter.scala 41:16]
  wire [3:0] _GEN_11 = 2'h1 == io_chosen ? io_in_1_bits_cmd : io_in_0_bits_cmd; // @[Arbiter.scala 41:16]
  wire [7:0] _GEN_12 = 2'h1 == io_chosen ? 8'hff : io_in_0_bits_wmask; // @[Arbiter.scala 41:16]
  wire [63:0] _GEN_13 = 2'h1 == io_chosen ? io_in_1_bits_wdata : io_in_0_bits_wdata; // @[Arbiter.scala 41:16]
  wire  _GEN_15 = 2'h2 == io_chosen ? io_in_2_valid : _GEN_8; // @[Arbiter.scala 41:16]
  wire [31:0] _GEN_16 = 2'h2 == io_chosen ? io_in_2_bits_addr : _GEN_9; // @[Arbiter.scala 41:16]
  wire [2:0] _GEN_17 = 2'h2 == io_chosen ? 3'h3 : _GEN_10; // @[Arbiter.scala 41:16]
  wire [3:0] _GEN_18 = 2'h2 == io_chosen ? io_in_2_bits_cmd : _GEN_11; // @[Arbiter.scala 41:16]
  wire [7:0] _GEN_19 = 2'h2 == io_chosen ? 8'hff : _GEN_12; // @[Arbiter.scala 41:16]
  wire [63:0] _GEN_20 = 2'h2 == io_chosen ? io_in_2_bits_wdata : _GEN_13; // @[Arbiter.scala 41:16]
  reg [2:0] value; // @[Counter.scala 29:33]
  reg [1:0] _T; // @[Arbiter.scala 46:22]
  wire  _T_1 = value != 3'h0; // @[Arbiter.scala 47:34]
  wire  _T_4 = io_out_bits_cmd[0] & io_out_bits_cmd[1]; // @[Crossbar.scala 100:62]
  wire  _T_5 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_6 = _T_5 & _T_4; // @[Arbiter.scala 50:25]
  wire [2:0] _T_9 = value + 3'h1; // @[Counter.scala 39:22]
  wire [1:0] _GEN_31 = io_in_2_valid ? 2'h2 : 2'h3; // @[Arbiter.scala 88:27]
  wire [1:0] _GEN_32 = io_in_1_valid ? 2'h1 : _GEN_31; // @[Arbiter.scala 88:27]
  wire [1:0] choice = io_in_0_valid ? 2'h0 : _GEN_32; // @[Arbiter.scala 88:27]
  wire  _T_10 = io_in_0_valid | io_in_1_valid; // @[Arbiter.scala 31:68]
  wire  _T_11 = _T_10 | io_in_2_valid; // @[Arbiter.scala 31:68]
  wire  _T_12 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  wire  _T_13 = ~_T_10; // @[Arbiter.scala 31:78]
  wire  _T_14 = ~_T_11; // @[Arbiter.scala 31:78]
  wire  _T_15 = _T == 2'h0; // @[Arbiter.scala 57:39]
  wire  _T_16 = _T_1 ? _T_15 : 1'h1; // @[Arbiter.scala 57:22]
  wire  _T_18 = _T == 2'h1; // @[Arbiter.scala 57:39]
  wire  _T_19 = _T_1 ? _T_18 : _T_12; // @[Arbiter.scala 57:22]
  wire  _T_21 = _T == 2'h2; // @[Arbiter.scala 57:39]
  wire  _T_22 = _T_1 ? _T_21 : _T_13; // @[Arbiter.scala 57:22]
  wire  _T_24 = _T == 2'h3; // @[Arbiter.scala 57:39]
  wire  _T_25 = _T_1 ? _T_24 : _T_14; // @[Arbiter.scala 57:22]
  assign io_in_0_ready = _T_16 & io_out_ready; // @[Arbiter.scala 57:16]
  assign io_in_1_ready = _T_19 & io_out_ready; // @[Arbiter.scala 57:16]
  assign io_in_2_ready = _T_22 & io_out_ready; // @[Arbiter.scala 57:16]
  assign io_in_3_ready = _T_25 & io_out_ready; // @[Arbiter.scala 57:16]
  assign io_out_valid = 2'h3 == io_chosen ? io_in_3_valid : _GEN_15; // @[Arbiter.scala 41:16]
  assign io_out_bits_addr = 2'h3 == io_chosen ? io_in_3_bits_addr : _GEN_16; // @[Arbiter.scala 42:15]
  assign io_out_bits_size = 2'h3 == io_chosen ? io_in_3_bits_size : _GEN_17; // @[Arbiter.scala 42:15]
  assign io_out_bits_cmd = 2'h3 == io_chosen ? io_in_3_bits_cmd : _GEN_18; // @[Arbiter.scala 42:15]
  assign io_out_bits_wmask = 2'h3 == io_chosen ? io_in_3_bits_wmask : _GEN_19; // @[Arbiter.scala 42:15]
  assign io_out_bits_wdata = 2'h3 == io_chosen ? io_in_3_bits_wdata : _GEN_20; // @[Arbiter.scala 42:15]
  assign io_chosen = _T_1 ? _T : choice; // @[Arbiter.scala 40:13 Arbiter.scala 55:31]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  _T = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 3'h0;
    end else if (_T_6) begin
      value <= _T_9;
    end
    if (_T_6) begin
      _T <= io_chosen;
    end
  end
endmodule
module SimpleBusCrossbarNto1_1(
  input         clock,
  input         reset,
  output        io_in_0_req_ready,
  input         io_in_0_req_valid,
  input  [31:0] io_in_0_req_bits_addr,
  input  [2:0]  io_in_0_req_bits_size,
  input  [3:0]  io_in_0_req_bits_cmd,
  input  [7:0]  io_in_0_req_bits_wmask,
  input  [63:0] io_in_0_req_bits_wdata,
  output        io_in_0_resp_valid,
  output [3:0]  io_in_0_resp_bits_cmd,
  output [63:0] io_in_0_resp_bits_rdata,
  output        io_in_1_req_ready,
  input         io_in_1_req_valid,
  input  [31:0] io_in_1_req_bits_addr,
  input  [3:0]  io_in_1_req_bits_cmd,
  input  [63:0] io_in_1_req_bits_wdata,
  output        io_in_1_resp_valid,
  output [3:0]  io_in_1_resp_bits_cmd,
  output [63:0] io_in_1_resp_bits_rdata,
  output        io_in_2_req_ready,
  input         io_in_2_req_valid,
  input  [31:0] io_in_2_req_bits_addr,
  input  [3:0]  io_in_2_req_bits_cmd,
  input  [63:0] io_in_2_req_bits_wdata,
  output        io_in_2_resp_valid,
  output [3:0]  io_in_2_resp_bits_cmd,
  output [63:0] io_in_2_resp_bits_rdata,
  output        io_in_3_req_ready,
  input         io_in_3_req_valid,
  input  [31:0] io_in_3_req_bits_addr,
  input  [2:0]  io_in_3_req_bits_size,
  input  [3:0]  io_in_3_req_bits_cmd,
  input  [7:0]  io_in_3_req_bits_wmask,
  input  [63:0] io_in_3_req_bits_wdata,
  input         io_in_3_resp_ready,
  output        io_in_3_resp_valid,
  output [3:0]  io_in_3_resp_bits_cmd,
  output [63:0] io_in_3_resp_bits_rdata,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [2:0]  io_out_req_bits_size,
  output [3:0]  io_out_req_bits_cmd,
  output [7:0]  io_out_req_bits_wmask,
  output [63:0] io_out_req_bits_wdata,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [3:0]  io_out_resp_bits_cmd,
  input  [63:0] io_out_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  inputArb_clock; // @[Crossbar.scala 101:24]
  wire  inputArb_reset; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_0_ready; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_0_valid; // @[Crossbar.scala 101:24]
  wire [31:0] inputArb_io_in_0_bits_addr; // @[Crossbar.scala 101:24]
  wire [2:0] inputArb_io_in_0_bits_size; // @[Crossbar.scala 101:24]
  wire [3:0] inputArb_io_in_0_bits_cmd; // @[Crossbar.scala 101:24]
  wire [7:0] inputArb_io_in_0_bits_wmask; // @[Crossbar.scala 101:24]
  wire [63:0] inputArb_io_in_0_bits_wdata; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_1_ready; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_1_valid; // @[Crossbar.scala 101:24]
  wire [31:0] inputArb_io_in_1_bits_addr; // @[Crossbar.scala 101:24]
  wire [3:0] inputArb_io_in_1_bits_cmd; // @[Crossbar.scala 101:24]
  wire [63:0] inputArb_io_in_1_bits_wdata; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_2_ready; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_2_valid; // @[Crossbar.scala 101:24]
  wire [31:0] inputArb_io_in_2_bits_addr; // @[Crossbar.scala 101:24]
  wire [3:0] inputArb_io_in_2_bits_cmd; // @[Crossbar.scala 101:24]
  wire [63:0] inputArb_io_in_2_bits_wdata; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_3_ready; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_3_valid; // @[Crossbar.scala 101:24]
  wire [31:0] inputArb_io_in_3_bits_addr; // @[Crossbar.scala 101:24]
  wire [2:0] inputArb_io_in_3_bits_size; // @[Crossbar.scala 101:24]
  wire [3:0] inputArb_io_in_3_bits_cmd; // @[Crossbar.scala 101:24]
  wire [7:0] inputArb_io_in_3_bits_wmask; // @[Crossbar.scala 101:24]
  wire [63:0] inputArb_io_in_3_bits_wdata; // @[Crossbar.scala 101:24]
  wire  inputArb_io_out_ready; // @[Crossbar.scala 101:24]
  wire  inputArb_io_out_valid; // @[Crossbar.scala 101:24]
  wire [31:0] inputArb_io_out_bits_addr; // @[Crossbar.scala 101:24]
  wire [2:0] inputArb_io_out_bits_size; // @[Crossbar.scala 101:24]
  wire [3:0] inputArb_io_out_bits_cmd; // @[Crossbar.scala 101:24]
  wire [7:0] inputArb_io_out_bits_wmask; // @[Crossbar.scala 101:24]
  wire [63:0] inputArb_io_out_bits_wdata; // @[Crossbar.scala 101:24]
  wire [1:0] inputArb_io_chosen; // @[Crossbar.scala 101:24]
  reg [1:0] state; // @[Crossbar.scala 98:22]
  wire  _T_1 = ~inputArb_io_out_bits_cmd[0]; // @[SimpleBus.scala 73:18]
  wire  _T_3 = ~inputArb_io_out_bits_cmd[3]; // @[SimpleBus.scala 73:29]
  wire  _T_4 = _T_1 & _T_3; // @[SimpleBus.scala 73:26]
  wire  _T_5 = ~_T_4; // @[Crossbar.scala 104:29]
  wire  _T_6 = inputArb_io_out_valid & _T_5; // @[Crossbar.scala 104:26]
  wire  _T_9 = _T_6 & _T_1; // @[Crossbar.scala 104:52]
  wire  _T_10 = ~_T_9; // @[Crossbar.scala 104:10]
  wire  _T_12 = _T_10 | reset; // @[Crossbar.scala 104:9]
  wire  _T_13 = ~_T_12; // @[Crossbar.scala 104:9]
  reg [1:0] inflightSrc; // @[Crossbar.scala 105:24]
  wire  _T_14 = state == 2'h0; // @[Crossbar.scala 109:47]
  wire  _GEN_58 = 2'h0 == inflightSrc; // @[Crossbar.scala 115:13]
  wire  _GEN_59 = 2'h1 == inflightSrc; // @[Crossbar.scala 115:13]
  wire  _GEN_60 = 2'h2 == inflightSrc; // @[Crossbar.scala 115:13]
  wire  _GEN_61 = 2'h3 == inflightSrc; // @[Crossbar.scala 115:13]
  wire  _T_18 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_19 = inputArb_io_out_ready & inputArb_io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_25 = inputArb_io_out_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_26 = inputArb_io_out_bits_cmd == 4'h1; // @[SimpleBus.scala 77:29]
  wire  _T_27 = _T_25 | _T_26; // @[Crossbar.scala 124:47]
  wire  _T_28 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_29 = io_out_resp_ready & io_out_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_30 = io_out_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire  _T_31 = _T_29 & _T_30; // @[Crossbar.scala 127:48]
  wire  _T_32 = 2'h2 == state; // @[Conditional.scala 37:30]
  LockingArbiter_1 inputArb ( // @[Crossbar.scala 101:24]
    .clock(inputArb_clock),
    .reset(inputArb_reset),
    .io_in_0_ready(inputArb_io_in_0_ready),
    .io_in_0_valid(inputArb_io_in_0_valid),
    .io_in_0_bits_addr(inputArb_io_in_0_bits_addr),
    .io_in_0_bits_size(inputArb_io_in_0_bits_size),
    .io_in_0_bits_cmd(inputArb_io_in_0_bits_cmd),
    .io_in_0_bits_wmask(inputArb_io_in_0_bits_wmask),
    .io_in_0_bits_wdata(inputArb_io_in_0_bits_wdata),
    .io_in_1_ready(inputArb_io_in_1_ready),
    .io_in_1_valid(inputArb_io_in_1_valid),
    .io_in_1_bits_addr(inputArb_io_in_1_bits_addr),
    .io_in_1_bits_cmd(inputArb_io_in_1_bits_cmd),
    .io_in_1_bits_wdata(inputArb_io_in_1_bits_wdata),
    .io_in_2_ready(inputArb_io_in_2_ready),
    .io_in_2_valid(inputArb_io_in_2_valid),
    .io_in_2_bits_addr(inputArb_io_in_2_bits_addr),
    .io_in_2_bits_cmd(inputArb_io_in_2_bits_cmd),
    .io_in_2_bits_wdata(inputArb_io_in_2_bits_wdata),
    .io_in_3_ready(inputArb_io_in_3_ready),
    .io_in_3_valid(inputArb_io_in_3_valid),
    .io_in_3_bits_addr(inputArb_io_in_3_bits_addr),
    .io_in_3_bits_size(inputArb_io_in_3_bits_size),
    .io_in_3_bits_cmd(inputArb_io_in_3_bits_cmd),
    .io_in_3_bits_wmask(inputArb_io_in_3_bits_wmask),
    .io_in_3_bits_wdata(inputArb_io_in_3_bits_wdata),
    .io_out_ready(inputArb_io_out_ready),
    .io_out_valid(inputArb_io_out_valid),
    .io_out_bits_addr(inputArb_io_out_bits_addr),
    .io_out_bits_size(inputArb_io_out_bits_size),
    .io_out_bits_cmd(inputArb_io_out_bits_cmd),
    .io_out_bits_wmask(inputArb_io_out_bits_wmask),
    .io_out_bits_wdata(inputArb_io_out_bits_wdata),
    .io_chosen(inputArb_io_chosen)
  );
  assign io_in_0_req_ready = inputArb_io_in_0_ready; // @[Crossbar.scala 102:68]
  assign io_in_0_resp_valid = _GEN_58 & io_out_resp_valid; // @[Crossbar.scala 113:26 Crossbar.scala 115:13]
  assign io_in_0_resp_bits_cmd = io_out_resp_bits_cmd; // @[Crossbar.scala 112:25]
  assign io_in_0_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 112:25]
  assign io_in_1_req_ready = inputArb_io_in_1_ready; // @[Crossbar.scala 102:68]
  assign io_in_1_resp_valid = _GEN_59 & io_out_resp_valid; // @[Crossbar.scala 113:26 Crossbar.scala 115:13]
  assign io_in_1_resp_bits_cmd = io_out_resp_bits_cmd; // @[Crossbar.scala 112:25]
  assign io_in_1_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 112:25]
  assign io_in_2_req_ready = inputArb_io_in_2_ready; // @[Crossbar.scala 102:68]
  assign io_in_2_resp_valid = _GEN_60 & io_out_resp_valid; // @[Crossbar.scala 113:26 Crossbar.scala 115:13]
  assign io_in_2_resp_bits_cmd = io_out_resp_bits_cmd; // @[Crossbar.scala 112:25]
  assign io_in_2_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 112:25]
  assign io_in_3_req_ready = inputArb_io_in_3_ready; // @[Crossbar.scala 102:68]
  assign io_in_3_resp_valid = _GEN_61 & io_out_resp_valid; // @[Crossbar.scala 113:26 Crossbar.scala 115:13]
  assign io_in_3_resp_bits_cmd = io_out_resp_bits_cmd; // @[Crossbar.scala 112:25]
  assign io_in_3_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 112:25]
  assign io_out_req_valid = inputArb_io_out_valid & _T_14; // @[Crossbar.scala 109:20]
  assign io_out_req_bits_addr = inputArb_io_out_bits_addr; // @[Crossbar.scala 107:19]
  assign io_out_req_bits_size = inputArb_io_out_bits_size; // @[Crossbar.scala 107:19]
  assign io_out_req_bits_cmd = inputArb_io_out_bits_cmd; // @[Crossbar.scala 107:19]
  assign io_out_req_bits_wmask = inputArb_io_out_bits_wmask; // @[Crossbar.scala 107:19]
  assign io_out_req_bits_wdata = inputArb_io_out_bits_wdata; // @[Crossbar.scala 107:19]
  assign io_out_resp_ready = 2'h3 == inflightSrc ? io_in_3_resp_ready : 1'h1; // @[Crossbar.scala 116:13]
  assign inputArb_clock = clock;
  assign inputArb_reset = reset;
  assign inputArb_io_in_0_valid = io_in_0_req_valid; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_addr = io_in_0_req_bits_addr; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_size = io_in_0_req_bits_size; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_cmd = io_in_0_req_bits_cmd; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_wmask = io_in_0_req_bits_wmask; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_wdata = io_in_0_req_bits_wdata; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_valid = io_in_1_req_valid; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_bits_addr = io_in_1_req_bits_addr; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_bits_cmd = io_in_1_req_bits_cmd; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_bits_wdata = io_in_1_req_bits_wdata; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_2_valid = io_in_2_req_valid; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_2_bits_addr = io_in_2_req_bits_addr; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_2_bits_cmd = io_in_2_req_bits_cmd; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_2_bits_wdata = io_in_2_req_bits_wdata; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_3_valid = io_in_3_req_valid; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_3_bits_addr = io_in_3_req_bits_addr; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_3_bits_size = io_in_3_req_bits_size; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_3_bits_cmd = io_in_3_req_bits_cmd; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_3_bits_wmask = io_in_3_req_bits_wmask; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_3_bits_wdata = io_in_3_req_bits_wdata; // @[Crossbar.scala 102:68]
  assign inputArb_io_out_ready = io_out_req_ready & _T_14; // @[Crossbar.scala 110:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  inflightSrc = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else if (_T_18) begin
      if (_T_19) begin
        if (_T_4) begin
          state <= 2'h1;
        end else if (_T_27) begin
          state <= 2'h2;
        end
      end
    end else if (_T_28) begin
      if (_T_31) begin
        state <= 2'h0;
      end
    end else if (_T_32) begin
      if (_T_29) begin
        state <= 2'h0;
      end
    end
    if (_T_18) begin
      if (_T_19) begin
        inflightSrc <= inputArb_io_chosen;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Crossbar.scala:104 assert(!(thisReq.valid && !thisReq.bits.isRead() && !thisReq.bits.isWrite()))\n"); // @[Crossbar.scala 104:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_13) begin
          $fatal; // @[Crossbar.scala 104:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module EmbeddedTLBExec(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [38:0]  io_in_bits_addr,
  input  [86:0]  io_in_bits_user,
  input          io_out_ready,
  output         io_out_valid,
  output [31:0]  io_out_bits_addr,
  output [86:0]  io_out_bits_user,
  input  [120:0] io_md_0,
  input  [120:0] io_md_1,
  input  [120:0] io_md_2,
  input  [120:0] io_md_3,
  output         io_mdWrite_wen,
  output         io_mdWrite_windex,
  output [3:0]   io_mdWrite_waymask,
  output [120:0] io_mdWrite_wdata,
  input          io_mdReady,
  input          io_mem_req_ready,
  output         io_mem_req_valid,
  output [31:0]  io_mem_req_bits_addr,
  output [2:0]   io_mem_req_bits_size,
  output [3:0]   io_mem_req_bits_cmd,
  output [7:0]   io_mem_req_bits_wmask,
  output [63:0]  io_mem_req_bits_wdata,
  output         io_mem_resp_ready,
  input          io_mem_resp_valid,
  input  [3:0]   io_mem_resp_bits_cmd,
  input  [63:0]  io_mem_resp_bits_rdata,
  input          io_flush,
  input  [63:0]  io_satp,
  input  [1:0]   io_pf_priviledgeMode,
  output         io_pf_loadPF,
  output         io_pf_storePF,
  output         io_ipf,
  output         io_isFinish,
  input          DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
`endif // RANDOMIZE_REG_INIT
  wire [8:0] vpn_vpn0 = io_in_bits_addr[20:12]; // @[EmbeddedTLB.scala 193:54]
  wire [8:0] vpn_vpn1 = io_in_bits_addr[29:21]; // @[EmbeddedTLB.scala 193:54]
  wire [8:0] vpn_vpn2 = io_in_bits_addr[38:30]; // @[EmbeddedTLB.scala 193:54]
  wire [19:0] satp_ppn = io_satp[19:0]; // @[EmbeddedTLB.scala 195:30]
  wire [15:0] satp_asid = io_satp[59:44]; // @[EmbeddedTLB.scala 195:30]
  wire  _T_39 = io_md_0[93:78] == satp_asid; // @[EmbeddedTLB.scala 204:117]
  wire  _T_40 = io_md_0[52] & _T_39; // @[EmbeddedTLB.scala 204:86]
  wire [17:0] _T_57 = {vpn_vpn2,vpn_vpn1}; // @[EmbeddedTLB.scala 204:201]
  wire [26:0] _T_58 = {vpn_vpn2,vpn_vpn1,vpn_vpn0}; // @[EmbeddedTLB.scala 204:201]
  wire [26:0] _T_59 = {9'h1ff,io_md_0[77:60]}; // @[Cat.scala 29:58]
  wire [26:0] _T_60 = _T_59 & io_md_0[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_62 = _T_59 & _T_58; // @[TLB.scala 131:84]
  wire  _T_63 = _T_60 == _T_62; // @[TLB.scala 131:48]
  wire  _T_64 = _T_40 & _T_63; // @[EmbeddedTLB.scala 204:132]
  wire  _T_91 = io_md_1[93:78] == satp_asid; // @[EmbeddedTLB.scala 204:117]
  wire  _T_92 = io_md_1[52] & _T_91; // @[EmbeddedTLB.scala 204:86]
  wire [26:0] _T_111 = {9'h1ff,io_md_1[77:60]}; // @[Cat.scala 29:58]
  wire [26:0] _T_112 = _T_111 & io_md_1[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_114 = _T_111 & _T_58; // @[TLB.scala 131:84]
  wire  _T_115 = _T_112 == _T_114; // @[TLB.scala 131:48]
  wire  _T_116 = _T_92 & _T_115; // @[EmbeddedTLB.scala 204:132]
  wire  _T_143 = io_md_2[93:78] == satp_asid; // @[EmbeddedTLB.scala 204:117]
  wire  _T_144 = io_md_2[52] & _T_143; // @[EmbeddedTLB.scala 204:86]
  wire [26:0] _T_163 = {9'h1ff,io_md_2[77:60]}; // @[Cat.scala 29:58]
  wire [26:0] _T_164 = _T_163 & io_md_2[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_166 = _T_163 & _T_58; // @[TLB.scala 131:84]
  wire  _T_167 = _T_164 == _T_166; // @[TLB.scala 131:48]
  wire  _T_168 = _T_144 & _T_167; // @[EmbeddedTLB.scala 204:132]
  wire  _T_195 = io_md_3[93:78] == satp_asid; // @[EmbeddedTLB.scala 204:117]
  wire  _T_196 = io_md_3[52] & _T_195; // @[EmbeddedTLB.scala 204:86]
  wire [26:0] _T_215 = {9'h1ff,io_md_3[77:60]}; // @[Cat.scala 29:58]
  wire [26:0] _T_216 = _T_215 & io_md_3[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_218 = _T_215 & _T_58; // @[TLB.scala 131:84]
  wire  _T_219 = _T_216 == _T_218; // @[TLB.scala 131:48]
  wire  _T_220 = _T_196 & _T_219; // @[EmbeddedTLB.scala 204:132]
  wire [3:0] hitVec = {_T_220,_T_168,_T_116,_T_64}; // @[EmbeddedTLB.scala 204:211]
  wire  _T_224 = |hitVec; // @[EmbeddedTLB.scala 205:35]
  wire  hit = io_in_valid & _T_224; // @[EmbeddedTLB.scala 205:25]
  wire  _T_226 = ~_T_224; // @[EmbeddedTLB.scala 206:29]
  wire  miss = io_in_valid & _T_226; // @[EmbeddedTLB.scala 206:26]
  reg [63:0] _T_227; // @[LFSR64.scala 25:23]
  wire  _T_230 = _T_227[0] ^ _T_227[1]; // @[LFSR64.scala 26:23]
  wire  _T_232 = _T_230 ^ _T_227[3]; // @[LFSR64.scala 26:33]
  wire  _T_234 = _T_232 ^ _T_227[4]; // @[LFSR64.scala 26:43]
  wire  _T_235 = _T_227 == 64'h0; // @[LFSR64.scala 28:24]
  wire [63:0] _T_237 = {_T_234,_T_227[63:1]}; // @[Cat.scala 29:58]
  wire [3:0] victimWaymask = 4'h1 << _T_227[1:0]; // @[EmbeddedTLB.scala 208:42]
  wire [3:0] waymask = hit ? hitVec : victimWaymask; // @[EmbeddedTLB.scala 209:20]
  wire [120:0] _T_244 = waymask[0] ? io_md_0 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_245 = waymask[1] ? io_md_1 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_246 = waymask[2] ? io_md_2 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_247 = waymask[3] ? io_md_3 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_248 = _T_244 | _T_245; // @[Mux.scala 27:72]
  wire [120:0] _T_249 = _T_248 | _T_246; // @[Mux.scala 27:72]
  wire [120:0] _T_250 = _T_249 | _T_247; // @[Mux.scala 27:72]
  wire [7:0] hitMeta_flag = _T_250[59:52]; // @[EmbeddedTLB.scala 215:70]
  wire [17:0] hitMeta_mask = _T_250[77:60]; // @[EmbeddedTLB.scala 215:70]
  wire [15:0] hitMeta_asid = _T_250[93:78]; // @[EmbeddedTLB.scala 215:70]
  wire [26:0] hitMeta_vpn = _T_250[120:94]; // @[EmbeddedTLB.scala 215:70]
  wire [31:0] hitData_pteaddr = _T_250[31:0]; // @[EmbeddedTLB.scala 216:70]
  wire [19:0] hitData_ppn = _T_250[51:32]; // @[EmbeddedTLB.scala 216:70]
  wire  hitFlag_v = hitMeta_flag[0]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_r = hitMeta_flag[1]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_w = hitMeta_flag[2]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_x = hitMeta_flag[3]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_u = hitMeta_flag[4]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_g = hitMeta_flag[5]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_a = hitMeta_flag[6]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_d = hitMeta_flag[7]; // @[EmbeddedTLB.scala 217:38]
  wire  _T_289 = ~hitFlag_a; // @[EmbeddedTLB.scala 221:23]
  wire  _T_294 = hit & _T_289; // @[EmbeddedTLB.scala 221:19]
  wire  _T_314 = io_pf_priviledgeMode == 2'h0; // @[EmbeddedTLB.scala 226:62]
  wire  _T_315 = ~hitFlag_u; // @[EmbeddedTLB.scala 226:75]
  wire  _T_316 = _T_314 & _T_315; // @[EmbeddedTLB.scala 226:72]
  wire  _T_317 = ~_T_316; // @[EmbeddedTLB.scala 226:42]
  wire  _T_318 = hit & _T_317; // @[EmbeddedTLB.scala 226:39]
  wire  _T_319 = io_pf_priviledgeMode == 2'h1; // @[EmbeddedTLB.scala 226:110]
  wire  _T_320 = _T_319 & hitFlag_u; // @[EmbeddedTLB.scala 226:120]
  wire  _T_324 = ~_T_320; // @[EmbeddedTLB.scala 226:90]
  wire  hitCheck = _T_318 & _T_324; // @[EmbeddedTLB.scala 226:87]
  wire  hitExec = hitCheck & hitFlag_x; // @[EmbeddedTLB.scala 227:26]
  wire  _T_329 = ~hitExec; // @[EmbeddedTLB.scala 239:42]
  wire  hitinstrPF = _T_329 & hit; // @[EmbeddedTLB.scala 239:52]
  wire  _T_295 = ~hitinstrPF; // @[EmbeddedTLB.scala 221:69]
  wire  _T_296 = _T_294 & _T_295; // @[EmbeddedTLB.scala 221:66]
  wire  _T_298 = io_pf_loadPF | io_pf_storePF; // @[Bundle.scala 135:23]
  wire  _T_300 = ~_T_298; // @[EmbeddedTLB.scala 221:84]
  wire  hitWB = _T_296 & _T_300; // @[EmbeddedTLB.scala 221:81]
  wire [7:0] _T_310 = {hitFlag_d,hitFlag_a,hitFlag_g,hitFlag_u,hitFlag_x,hitFlag_w,hitFlag_r,hitFlag_v}; // @[EmbeddedTLB.scala 222:79]
  wire [7:0] hitRefillFlag = 8'h40 | _T_310; // @[EmbeddedTLB.scala 222:69]
  wire [39:0] _T_313 = {10'h0,hitData_ppn,2'h0,hitRefillFlag}; // @[Cat.scala 29:58]
  reg [39:0] hitWBStore; // @[Reg.scala 15:16]
  wire  hitLoad = hitCheck & hitFlag_r; // @[EmbeddedTLB.scala 228:26]
  wire  hitStore = hitCheck & hitFlag_w; // @[EmbeddedTLB.scala 229:27]
  reg [2:0] state; // @[EmbeddedTLB.scala 247:22]
  reg [1:0] level; // @[EmbeddedTLB.scala 248:22]
  reg [63:0] memRespStore; // @[EmbeddedTLB.scala 250:25]
  reg [17:0] missMaskStore; // @[EmbeddedTLB.scala 252:26]
  wire  memRdata_flag_v = io_mem_resp_bits_rdata[0]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_r = io_mem_resp_bits_rdata[1]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_w = io_mem_resp_bits_rdata[2]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_x = io_mem_resp_bits_rdata[3]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_u = io_mem_resp_bits_rdata[4]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_g = io_mem_resp_bits_rdata[5]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_a = io_mem_resp_bits_rdata[6]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_d = io_mem_resp_bits_rdata[7]; // @[EmbeddedTLB.scala 255:49]
  wire [1:0] memRdata_rsw = io_mem_resp_bits_rdata[9:8]; // @[EmbeddedTLB.scala 255:49]
  wire [19:0] memRdata_ppn = io_mem_resp_bits_rdata[29:10]; // @[EmbeddedTLB.scala 255:49]
  wire [33:0] memRdata_reserved = io_mem_resp_bits_rdata[63:30]; // @[EmbeddedTLB.scala 255:49]
  reg [31:0] raddr; // @[EmbeddedTLB.scala 256:18]
  wire  _T_343 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  reg  alreadyOutFire; // @[Reg.scala 27:20]
  wire  _GEN_2 = _T_343 | alreadyOutFire; // @[Reg.scala 28:19]
  reg  needFlush; // @[EmbeddedTLB.scala 260:26]
  wire  isFlush = needFlush | io_flush; // @[EmbeddedTLB.scala 262:27]
  wire  _T_344 = state != 3'h0; // @[EmbeddedTLB.scala 263:27]
  wire  _T_345 = io_flush & _T_344; // @[EmbeddedTLB.scala 263:17]
  wire  _GEN_3 = _T_345 | needFlush; // @[EmbeddedTLB.scala 263:40]
  wire  _T_347 = _T_343 & needFlush; // @[EmbeddedTLB.scala 264:23]
  wire  _GEN_4 = _T_347 ? 1'h0 : _GEN_3; // @[EmbeddedTLB.scala 264:37]
  reg  missIPF; // @[EmbeddedTLB.scala 266:24]
  wire  _T_348 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_349 = ~io_flush; // @[EmbeddedTLB.scala 271:13]
  wire  _T_350 = _T_349 & hitWB; // @[EmbeddedTLB.scala 271:22]
  wire  _T_352 = miss & _T_349; // @[EmbeddedTLB.scala 275:24]
  wire [31:0] _T_354 = {satp_ppn,vpn_vpn2,3'h0}; // @[Cat.scala 29:58]
  wire  _T_355 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_356 = io_mem_req_ready & io_mem_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_357 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire [7:0] _T_365 = {memRdata_flag_d,memRdata_flag_a,memRdata_flag_g,memRdata_flag_u,memRdata_flag_x,memRdata_flag_w,memRdata_flag_r,memRdata_flag_v}; // @[EmbeddedTLB.scala 292:44]
  wire  _T_375 = io_mem_resp_ready & io_mem_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_376 = _T_365[1] | _T_365[3]; // @[EmbeddedTLB.scala 297:34]
  wire  _T_377 = ~_T_376; // @[EmbeddedTLB.scala 297:21]
  wire  _T_378 = level == 2'h3; // @[EmbeddedTLB.scala 297:58]
  wire  _T_379 = level == 2'h2; // @[EmbeddedTLB.scala 297:73]
  wire  _T_380 = _T_378 | _T_379; // @[EmbeddedTLB.scala 297:65]
  wire  _T_381 = _T_377 & _T_380; // @[EmbeddedTLB.scala 297:49]
  wire  _T_382 = ~_T_365[0]; // @[EmbeddedTLB.scala 298:16]
  wire  _T_383 = ~_T_365[1]; // @[EmbeddedTLB.scala 298:32]
  wire  _T_384 = _T_383 & _T_365[2]; // @[EmbeddedTLB.scala 298:44]
  wire  _T_385 = _T_382 | _T_384; // @[EmbeddedTLB.scala 298:28]
  reg [63:0] _T_386; // @[GTimer.scala 24:20]
  wire [63:0] _T_388 = _T_386 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_392 = ~reset; // @[Debug.scala 56:24]
  wire [8:0] _T_417 = _T_378 ? vpn_vpn1 : vpn_vpn0; // @[EmbeddedTLB.scala 311:50]
  wire [31:0] _T_419 = {memRdata_ppn,_T_417,3'h0}; // @[Cat.scala 29:58]
  wire  _GEN_19 = _T_385 | missIPF; // @[EmbeddedTLB.scala 298:60]
  wire  _T_420 = level != 2'h0; // @[EmbeddedTLB.scala 313:27]
  wire  _T_422 = ~_T_365[4]; // @[EmbeddedTLB.scala 314:74]
  wire  _T_423 = _T_314 & _T_422; // @[EmbeddedTLB.scala 314:71]
  wire  _T_424 = ~_T_423; // @[EmbeddedTLB.scala 314:41]
  wire  _T_425 = _T_365[0] & _T_424; // @[EmbeddedTLB.scala 314:38]
  wire  _T_427 = _T_319 & _T_365[4]; // @[EmbeddedTLB.scala 314:120]
  wire  _T_431 = ~_T_427; // @[EmbeddedTLB.scala 314:90]
  wire  _T_432 = _T_425 & _T_431; // @[EmbeddedTLB.scala 314:87]
  wire  _T_433 = _T_432 & _T_365[3]; // @[EmbeddedTLB.scala 315:36]
  wire [7:0] _T_451 = {_T_365[7],_T_365[6],_T_365[5],_T_365[4],_T_365[3],_T_365[2],_T_365[1],_T_365[0]}; // @[EmbeddedTLB.scala 320:79]
  wire [7:0] _T_452 = 8'h40 | _T_451; // @[EmbeddedTLB.scala 320:68]
  wire [63:0] _T_453 = io_mem_resp_bits_rdata | 64'h40; // @[EmbeddedTLB.scala 321:50]
  wire  _T_454 = ~_T_433; // @[EmbeddedTLB.scala 323:19]
  wire  _GEN_21 = _T_454 | missIPF; // @[EmbeddedTLB.scala 323:30]
  wire  _GEN_23 = _T_454 ? 1'h0 : 1'h1; // @[EmbeddedTLB.scala 323:30]
  wire [17:0] _T_458 = _T_379 ? 18'h3fe00 : 18'h3ffff; // @[EmbeddedTLB.scala 339:59]
  wire [17:0] _T_459 = _T_378 ? 18'h0 : _T_458; // @[EmbeddedTLB.scala 339:26]
  wire [7:0] _GEN_24 = _T_420 ? _T_452 : 8'h0; // @[EmbeddedTLB.scala 313:36]
  wire  _GEN_28 = _T_420 & _GEN_23; // @[EmbeddedTLB.scala 313:36]
  wire [17:0] _GEN_29 = _T_420 ? _T_459 : 18'h3ffff; // @[EmbeddedTLB.scala 313:36]
  wire [17:0] _GEN_37 = _T_381 ? 18'h3ffff : _GEN_29; // @[EmbeddedTLB.scala 297:82]
  wire [17:0] _GEN_45 = isFlush ? 18'h3ffff : _GEN_37; // @[EmbeddedTLB.scala 294:24]
  wire [17:0] _GEN_54 = _T_375 ? _GEN_45 : 18'h3ffff; // @[EmbeddedTLB.scala 293:33]
  wire [17:0] _GEN_77 = _T_357 ? _GEN_54 : 18'h3ffff; // @[Conditional.scala 39:67]
  wire [17:0] _GEN_88 = _T_355 ? 18'h3ffff : _GEN_77; // @[Conditional.scala 39:67]
  wire [17:0] missMask = _T_348 ? 18'h3ffff : _GEN_88; // @[Conditional.scala 40:58]
  wire [7:0] _GEN_34 = _T_381 ? 8'h0 : _GEN_24; // @[EmbeddedTLB.scala 297:82]
  wire  _GEN_36 = _T_381 ? 1'h0 : _GEN_28; // @[EmbeddedTLB.scala 297:82]
  wire [7:0] _GEN_42 = isFlush ? 8'h0 : _GEN_34; // @[EmbeddedTLB.scala 294:24]
  wire  _GEN_44 = isFlush ? 1'h0 : _GEN_36; // @[EmbeddedTLB.scala 294:24]
  wire [1:0] _T_461 = level - 2'h1; // @[EmbeddedTLB.scala 342:24]
  wire [7:0] _GEN_51 = _T_375 ? _GEN_42 : 8'h0; // @[EmbeddedTLB.scala 293:33]
  wire  _GEN_53 = _T_375 & _GEN_44; // @[EmbeddedTLB.scala 293:33]
  wire  _T_462 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_464 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_466 = _T_343 | io_flush; // @[EmbeddedTLB.scala 353:44]
  wire  _T_467 = _T_466 | alreadyOutFire; // @[EmbeddedTLB.scala 353:55]
  wire  _T_468 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire [7:0] _GEN_74 = _T_357 ? _GEN_51 : 8'h0; // @[Conditional.scala 39:67]
  wire  _GEN_76 = _T_357 & _GEN_53; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_85 = _T_355 ? 8'h0 : _GEN_74; // @[Conditional.scala 39:67]
  wire  _GEN_87 = _T_355 ? 1'h0 : _GEN_76; // @[Conditional.scala 39:67]
  wire [7:0] missRefillFlag = _T_348 ? 8'h0 : _GEN_85; // @[Conditional.scala 40:58]
  wire  missMetaRefill = _T_348 ? 1'h0 : _GEN_87; // @[Conditional.scala 40:58]
  wire  cmd = state == 3'h3; // @[EmbeddedTLB.scala 365:23]
  wire  _T_472 = state == 3'h1; // @[EmbeddedTLB.scala 367:31]
  wire  _T_474 = _T_472 | cmd; // @[EmbeddedTLB.scala 367:48]
  wire  _T_475 = ~isFlush; // @[EmbeddedTLB.scala 367:77]
  wire  _T_478 = missMetaRefill & _T_475; // @[EmbeddedTLB.scala 371:50]
  wire  _T_479 = state == 3'h0; // @[EmbeddedTLB.scala 371:82]
  wire  _T_480 = hitWB & _T_479; // @[EmbeddedTLB.scala 371:73]
  wire  _T_482 = _T_480 & _T_475; // @[EmbeddedTLB.scala 371:93]
  wire  _T_483 = _T_478 | _T_482; // @[EmbeddedTLB.scala 371:63]
  reg  _T_484; // @[EmbeddedTLB.scala 371:33]
  reg  _T_490; // @[EmbeddedTLB.scala 372:21]
  reg [3:0] _T_491; // @[EmbeddedTLB.scala 372:60]
  reg [26:0] _T_494; // @[EmbeddedTLB.scala 372:84]
  reg [15:0] _T_496; // @[EmbeddedTLB.scala 373:19]
  reg [17:0] _T_498; // @[EmbeddedTLB.scala 373:72]
  reg [7:0] _T_500; // @[EmbeddedTLB.scala 374:19]
  reg [19:0] _T_502; // @[EmbeddedTLB.scala 374:77]
  reg [31:0] _T_504; // @[EmbeddedTLB.scala 375:22]
  wire [59:0] _T_506 = {_T_500,_T_502,_T_504}; // @[Cat.scala 29:58]
  wire [60:0] _T_508 = {_T_494,_T_496,_T_498}; // @[Cat.scala 29:58]
  wire [31:0] _T_511 = {hitData_ppn,12'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_514 = {2'h3,hitMeta_mask,12'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_515 = _T_511 & _T_514; // @[BitUtils.scala 32:13]
  wire [31:0] _T_516 = ~_T_514; // @[BitUtils.scala 32:38]
  wire [31:0] _T_517 = io_in_bits_addr[31:0] & _T_516; // @[BitUtils.scala 32:36]
  wire [31:0] _T_518 = _T_515 | _T_517; // @[BitUtils.scala 32:25]
  wire [31:0] _T_533 = {memRespStore[29:10],12'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_536 = {2'h3,missMaskStore,12'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_537 = _T_533 & _T_536; // @[BitUtils.scala 32:13]
  wire [31:0] _T_538 = ~_T_536; // @[BitUtils.scala 32:38]
  wire [31:0] _T_539 = io_in_bits_addr[31:0] & _T_538; // @[BitUtils.scala 32:36]
  wire [31:0] _T_540 = _T_537 | _T_539; // @[BitUtils.scala 32:25]
  wire  _T_542 = ~hitWB; // @[EmbeddedTLB.scala 380:45]
  wire  _T_543 = hit & _T_542; // @[EmbeddedTLB.scala 380:42]
  wire  _T_548 = state == 3'h4; // @[EmbeddedTLB.scala 380:97]
  wire  _T_549 = _T_543 ? _T_300 : _T_548; // @[EmbeddedTLB.scala 380:37]
  wire  _T_552 = io_out_ready & _T_479; // @[EmbeddedTLB.scala 382:31]
  wire  _T_553 = ~miss; // @[EmbeddedTLB.scala 382:56]
  wire  _T_554 = _T_552 & _T_553; // @[EmbeddedTLB.scala 382:53]
  wire  _T_556 = _T_554 & _T_542; // @[EmbeddedTLB.scala 382:62]
  wire  _T_557 = _T_556 & io_mdReady; // @[EmbeddedTLB.scala 382:72]
  reg [63:0] _T_569; // @[GTimer.scala 24:20]
  wire [63:0] _T_571 = _T_569 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_578; // @[GTimer.scala 24:20]
  wire [63:0] _T_580 = _T_578 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_594; // @[GTimer.scala 24:20]
  wire [63:0] _T_596 = _T_594 + 64'h1; // @[GTimer.scala 25:12]
  wire [4:0] _T_606 = {memRdata_flag_u,memRdata_flag_x,memRdata_flag_w,memRdata_flag_r,memRdata_flag_v}; // @[EmbeddedTLB.scala 390:145]
  wire [63:0] _T_612 = {memRdata_reserved,memRdata_ppn,memRdata_rsw,memRdata_flag_d,memRdata_flag_a,memRdata_flag_g,_T_606}; // @[EmbeddedTLB.scala 390:145]
  reg [63:0] _T_613; // @[GTimer.scala 24:20]
  wire [63:0] _T_615 = _T_613 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_718; // @[GTimer.scala 24:20]
  wire [63:0] _T_720 = _T_718 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_783; // @[GTimer.scala 24:20]
  wire [63:0] _T_785 = _T_783 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_792; // @[GTimer.scala 24:20]
  wire [63:0] _T_794 = _T_792 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_801; // @[GTimer.scala 24:20]
  wire [63:0] _T_803 = _T_801 + 64'h1; // @[GTimer.scala 25:12]
  wire  _GEN_104 = ~_T_348; // @[Debug.scala 56:24]
  wire  _GEN_105 = ~_T_355; // @[Debug.scala 56:24]
  wire  _GEN_106 = _GEN_104 & _GEN_105; // @[Debug.scala 56:24]
  wire  _GEN_107 = _GEN_106 & _T_357; // @[Debug.scala 56:24]
  wire  _GEN_108 = _GEN_107 & _T_375; // @[Debug.scala 56:24]
  wire  _GEN_110 = _GEN_108 & _T_475; // @[Debug.scala 56:24]
  wire  _GEN_111 = _GEN_110 & _T_381; // @[Debug.scala 56:24]
  wire  _GEN_112 = _GEN_111 & _T_385; // @[Debug.scala 56:24]
  wire  _GEN_113 = _GEN_112 & DISPLAY_ENABLE; // @[Debug.scala 56:24]
  assign io_in_ready = _T_557 & _T_300; // @[EmbeddedTLB.scala 382:15]
  assign io_out_valid = io_in_valid & _T_549; // @[EmbeddedTLB.scala 380:16]
  assign io_out_bits_addr = hit ? _T_518 : _T_540; // @[EmbeddedTLB.scala 378:15 EmbeddedTLB.scala 379:20]
  assign io_out_bits_user = io_in_bits_user; // @[EmbeddedTLB.scala 378:15]
  assign io_mdWrite_wen = _T_484; // @[TLB.scala 214:14]
  assign io_mdWrite_windex = _T_490; // @[TLB.scala 215:17]
  assign io_mdWrite_waymask = _T_491; // @[TLB.scala 216:18]
  assign io_mdWrite_wdata = {_T_508,_T_506}; // @[TLB.scala 217:16]
  assign io_mem_req_valid = _T_474 & _T_475; // @[EmbeddedTLB.scala 367:20]
  assign io_mem_req_bits_addr = hitWB ? hitData_pteaddr : raddr; // @[SimpleBus.scala 64:15]
  assign io_mem_req_bits_size = 3'h3; // @[SimpleBus.scala 66:15]
  assign io_mem_req_bits_cmd = {{3'd0}, cmd}; // @[SimpleBus.scala 65:14]
  assign io_mem_req_bits_wmask = 8'hff; // @[SimpleBus.scala 68:16]
  assign io_mem_req_bits_wdata = hitWB ? {{24'd0}, hitWBStore} : memRespStore; // @[SimpleBus.scala 67:16]
  assign io_mem_resp_ready = 1'h1; // @[EmbeddedTLB.scala 368:21]
  assign io_pf_loadPF = 1'h0; // @[EmbeddedTLB.scala 199:13 EmbeddedTLB.scala 236:16]
  assign io_pf_storePF = 1'h0; // @[EmbeddedTLB.scala 200:14 EmbeddedTLB.scala 237:17]
  assign io_ipf = hit ? hitinstrPF : missIPF; // @[EmbeddedTLB.scala 384:10]
  assign io_isFinish = _T_343 | _T_298; // @[EmbeddedTLB.scala 385:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  _T_227 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  hitWBStore = _RAND_1[39:0];
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  level = _RAND_3[1:0];
  _RAND_4 = {2{`RANDOM}};
  memRespStore = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  missMaskStore = _RAND_5[17:0];
  _RAND_6 = {1{`RANDOM}};
  raddr = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  alreadyOutFire = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  needFlush = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  missIPF = _RAND_9[0:0];
  _RAND_10 = {2{`RANDOM}};
  _T_386 = _RAND_10[63:0];
  _RAND_11 = {1{`RANDOM}};
  _T_484 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _T_490 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _T_491 = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  _T_494 = _RAND_14[26:0];
  _RAND_15 = {1{`RANDOM}};
  _T_496 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  _T_498 = _RAND_16[17:0];
  _RAND_17 = {1{`RANDOM}};
  _T_500 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  _T_502 = _RAND_18[19:0];
  _RAND_19 = {1{`RANDOM}};
  _T_504 = _RAND_19[31:0];
  _RAND_20 = {2{`RANDOM}};
  _T_569 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  _T_578 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  _T_594 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  _T_613 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  _T_718 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  _T_783 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  _T_792 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  _T_801 = _RAND_27[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_227 <= 64'h1234567887654321;
    end else if (_T_235) begin
      _T_227 <= 64'h1;
    end else begin
      _T_227 <= _T_237;
    end
    if (hitWB) begin
      hitWBStore <= _T_313;
    end
    if (reset) begin
      state <= 3'h0;
    end else if (_T_348) begin
      if (_T_350) begin
        state <= 3'h3;
      end else if (_T_352) begin
        state <= 3'h1;
      end
    end else if (_T_355) begin
      if (isFlush) begin
        state <= 3'h0;
      end else if (_T_356) begin
        state <= 3'h2;
      end
    end else if (_T_357) begin
      if (_T_375) begin
        if (isFlush) begin
          state <= 3'h0;
        end else if (_T_381) begin
          if (_T_385) begin
            state <= 3'h4;
          end else begin
            state <= 3'h1;
          end
        end else if (_T_420) begin
          state <= 3'h4;
        end
      end
    end else if (_T_462) begin
      if (isFlush) begin
        state <= 3'h0;
      end else if (_T_356) begin
        state <= 3'h4;
      end
    end else if (_T_464) begin
      if (_T_467) begin
        state <= 3'h0;
      end
    end else if (_T_468) begin
      state <= 3'h0;
    end
    if (reset) begin
      level <= 2'h3;
    end else if (_T_348) begin
      if (!(_T_350)) begin
        if (_T_352) begin
          level <= 2'h3;
        end
      end
    end else if (!(_T_355)) begin
      if (_T_357) begin
        if (_T_375) begin
          level <= _T_461;
        end
      end
    end
    if (!(_T_348)) begin
      if (!(_T_355)) begin
        if (_T_357) begin
          if (_T_375) begin
            if (!(isFlush)) begin
              if (!(_T_381)) begin
                if (_T_420) begin
                  memRespStore <= _T_453;
                end
              end
            end
          end
        end
      end
    end
    if (!(_T_348)) begin
      if (!(_T_355)) begin
        if (_T_357) begin
          if (_T_375) begin
            if (!(isFlush)) begin
              if (!(_T_381)) begin
                if (_T_420) begin
                  if (_T_348) begin
                    missMaskStore <= 18'h3ffff;
                  end else if (_T_355) begin
                    missMaskStore <= 18'h3ffff;
                  end else if (_T_357) begin
                    if (_T_375) begin
                      if (isFlush) begin
                        missMaskStore <= 18'h3ffff;
                      end else if (_T_381) begin
                        missMaskStore <= 18'h3ffff;
                      end else if (_T_420) begin
                        if (_T_378) begin
                          missMaskStore <= 18'h0;
                        end else if (_T_379) begin
                          missMaskStore <= 18'h3fe00;
                        end else begin
                          missMaskStore <= 18'h3ffff;
                        end
                      end else begin
                        missMaskStore <= 18'h3ffff;
                      end
                    end else begin
                      missMaskStore <= 18'h3ffff;
                    end
                  end else begin
                    missMaskStore <= 18'h3ffff;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_348) begin
      if (!(_T_350)) begin
        if (_T_352) begin
          raddr <= _T_354;
        end
      end
    end else if (!(_T_355)) begin
      if (_T_357) begin
        if (_T_375) begin
          if (!(isFlush)) begin
            if (_T_381) begin
              if (!(_T_385)) begin
                raddr <= _T_419;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      alreadyOutFire <= 1'h0;
    end else if (_T_348) begin
      if (_T_350) begin
        alreadyOutFire <= 1'h0;
      end else if (_T_352) begin
        alreadyOutFire <= 1'h0;
      end else begin
        alreadyOutFire <= _GEN_2;
      end
    end else if (_T_355) begin
      alreadyOutFire <= _GEN_2;
    end else if (_T_357) begin
      alreadyOutFire <= _GEN_2;
    end else if (_T_462) begin
      alreadyOutFire <= _GEN_2;
    end else if (_T_464) begin
      if (_T_467) begin
        alreadyOutFire <= 1'h0;
      end else begin
        alreadyOutFire <= _GEN_2;
      end
    end else begin
      alreadyOutFire <= _GEN_2;
    end
    if (reset) begin
      needFlush <= 1'h0;
    end else if (_T_348) begin
      if (_T_350) begin
        needFlush <= 1'h0;
      end else if (_T_352) begin
        needFlush <= 1'h0;
      end else if (_T_347) begin
        needFlush <= 1'h0;
      end else begin
        needFlush <= _GEN_3;
      end
    end else if (_T_355) begin
      if (isFlush) begin
        needFlush <= 1'h0;
      end else if (_T_347) begin
        needFlush <= 1'h0;
      end else begin
        needFlush <= _GEN_3;
      end
    end else if (_T_357) begin
      if (_T_375) begin
        if (isFlush) begin
          needFlush <= 1'h0;
        end else if (_T_347) begin
          needFlush <= 1'h0;
        end else begin
          needFlush <= _GEN_3;
        end
      end else if (_T_347) begin
        needFlush <= 1'h0;
      end else begin
        needFlush <= _GEN_3;
      end
    end else if (_T_462) begin
      if (isFlush) begin
        needFlush <= 1'h0;
      end else begin
        needFlush <= _GEN_4;
      end
    end else begin
      needFlush <= _GEN_4;
    end
    if (reset) begin
      missIPF <= 1'h0;
    end else if (!(_T_348)) begin
      if (!(_T_355)) begin
        if (_T_357) begin
          if (_T_375) begin
            if (!(isFlush)) begin
              if (_T_381) begin
                missIPF <= _GEN_19;
              end else if (_T_420) begin
                missIPF <= _GEN_21;
              end
            end
          end
        end else if (!(_T_462)) begin
          if (_T_464) begin
            if (_T_467) begin
              missIPF <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_386 <= 64'h0;
    end else begin
      _T_386 <= _T_388;
    end
    if (reset) begin
      _T_484 <= 1'h0;
    end else begin
      _T_484 <= _T_483;
    end
    _T_490 <= io_in_bits_addr[12];
    if (hit) begin
      _T_491 <= hitVec;
    end else begin
      _T_491 <= victimWaymask;
    end
    _T_494 <= {_T_57,vpn_vpn0};
    if (hitWB) begin
      _T_496 <= hitMeta_asid;
    end else begin
      _T_496 <= satp_asid;
    end
    if (hitWB) begin
      _T_498 <= hitMeta_mask;
    end else if (_T_348) begin
      _T_498 <= 18'h3ffff;
    end else if (_T_355) begin
      _T_498 <= 18'h3ffff;
    end else if (_T_357) begin
      if (_T_375) begin
        if (isFlush) begin
          _T_498 <= 18'h3ffff;
        end else if (_T_381) begin
          _T_498 <= 18'h3ffff;
        end else if (_T_420) begin
          if (_T_378) begin
            _T_498 <= 18'h0;
          end else if (_T_379) begin
            _T_498 <= 18'h3fe00;
          end else begin
            _T_498 <= 18'h3ffff;
          end
        end else begin
          _T_498 <= 18'h3ffff;
        end
      end else begin
        _T_498 <= 18'h3ffff;
      end
    end else begin
      _T_498 <= 18'h3ffff;
    end
    if (hitWB) begin
      _T_500 <= hitRefillFlag;
    end else if (_T_348) begin
      _T_500 <= 8'h0;
    end else if (_T_355) begin
      _T_500 <= 8'h0;
    end else if (_T_357) begin
      if (_T_375) begin
        if (isFlush) begin
          _T_500 <= 8'h0;
        end else if (_T_381) begin
          _T_500 <= 8'h0;
        end else if (_T_420) begin
          _T_500 <= _T_452;
        end else begin
          _T_500 <= 8'h0;
        end
      end else begin
        _T_500 <= 8'h0;
      end
    end else begin
      _T_500 <= 8'h0;
    end
    if (hitWB) begin
      _T_502 <= hitData_ppn;
    end else begin
      _T_502 <= memRdata_ppn;
    end
    if (hitWB) begin
      _T_504 <= hitData_pteaddr;
    end else begin
      _T_504 <= raddr;
    end
    if (reset) begin
      _T_569 <= 64'h0;
    end else begin
      _T_569 <= _T_571;
    end
    if (reset) begin
      _T_578 <= 64'h0;
    end else begin
      _T_578 <= _T_580;
    end
    if (reset) begin
      _T_594 <= 64'h0;
    end else begin
      _T_594 <= _T_596;
    end
    if (reset) begin
      _T_613 <= 64'h0;
    end else begin
      _T_613 <= _T_615;
    end
    if (reset) begin
      _T_718 <= 64'h0;
    end else begin
      _T_718 <= _T_720;
    end
    if (reset) begin
      _T_783 <= 64'h0;
    end else begin
      _T_783 <= _T_785;
    end
    if (reset) begin
      _T_792 <= 64'h0;
    end else begin
      _T_792 <= _T_794;
    end
    if (reset) begin
      _T_801 <= 64'h0;
    end else begin
      _T_801 <= _T_803;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_113 & _T_392) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec: ",_T_386); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_113 & _T_392) begin
          $fwrite(32'h80000002,"tlbException!!! "); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_113 & _T_392) begin
          $fwrite(32'h80000002," req:addr = 0x%x, cmd = %d, size = %d, wmask = 0x%x, wdata = 0x%x  Memreq:DecoupledIO(ready -> %d, valid -> %d, bits -> addr = 0x%x, cmd = %d, size = %d, wmask = 0x%x, wdata = 0x%x)  MemResp:DecoupledIO(ready -> %d, valid -> %d, bits -> rdata = %x, cmd = %d)",io_in_bits_addr,4'h0,3'h3,8'h0,64'h0,io_mem_req_ready,io_mem_req_valid,io_mem_req_bits_addr,io_mem_req_bits_cmd,io_mem_req_bits_size,io_mem_req_bits_wmask,io_mem_req_bits_wdata,io_mem_resp_ready,io_mem_resp_valid,io_mem_resp_bits_rdata,io_mem_resp_bits_cmd); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_113 & _T_392) begin
          $fwrite(32'h80000002," level:%d",level); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_113 & _T_392) begin
          $fwrite(32'h80000002,"\n"); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_392) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec: ",_T_569); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_392) begin
          $fwrite(32'h80000002,"In(%d, %d) Out(%d, %d) InAddr:%x OutAddr:%x cmd:%d \n",io_in_valid,io_in_ready,io_out_valid,io_out_ready,io_in_bits_addr,io_out_bits_addr,4'h0); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_392) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec: ",_T_578); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_392) begin
          $fwrite(32'h80000002,"isAMO:%d io.Flush:%d needFlush:%d alreadyOutFire:%d isFinish:%d\n",1'h0,io_flush,needFlush,alreadyOutFire,io_isFinish); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_392) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec: ",_T_594); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_392) begin
          $fwrite(32'h80000002,"hit:%d hitWB:%d hitVPN:%x hitFlag:%x hitPPN:%x hitRefillFlag:%x hitWBStore:%x hitCheck:%d hitExec:%d hitLoad:%d hitStore:%d\n",hit,hitWB,hitMeta_vpn,_T_310,hitData_ppn,hitRefillFlag,hitWBStore,hitCheck,hitExec,hitLoad,hitStore); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_392) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec: ",_T_613); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_392) begin
          $fwrite(32'h80000002,"miss:%d state:%d level:%d raddr:%x memRdata:%x missMask:%x missRefillFlag:%x missMetaRefill:%d\n",miss,state,level,raddr,_T_612,missMask,missRefillFlag,missMetaRefill); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_392) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec: ",_T_718); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_392) begin
          $fwrite(32'h80000002,"meta/data: (0)%x|%b|%x (1)%x|%b|%x (2)%x|%b|%x (3)%x|%b|%x rread:%d\n",io_md_0[120:94],io_md_0[59:52],io_md_0[51:32],io_md_1[120:94],io_md_1[59:52],io_md_1[51:32],io_md_2[120:94],io_md_2[59:52],io_md_2[51:32],io_md_3[120:94],io_md_3[59:52],io_md_3[51:32],io_mdReady); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_392) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec: ",_T_783); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_392) begin
          $fwrite(32'h80000002,"md: wen:%d windex:%x waymask:%x vpn:%x asid:%x mask:%x flag:%x asid:%x ppn:%x pteaddr:%x\n",io_mdWrite_wen,io_mdWrite_windex,io_mdWrite_waymask,io_mdWrite_wdata[120:94],io_mdWrite_wdata[93:78],io_mdWrite_wdata[77:60],io_mdWrite_wdata[59:52],io_mdWrite_wdata[93:78],io_mdWrite_wdata[51:32],io_mdWrite_wdata[31:0]); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_392) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec: ",_T_792); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_392) begin
          $fwrite(32'h80000002,"MemReq(%d, %d) MemResp(%d, %d) addr:%x cmd:%d rdata:%x cmd:%d\n",io_mem_req_valid,io_mem_req_ready,io_mem_resp_valid,io_mem_resp_ready,io_mem_req_bits_addr,io_mem_req_bits_cmd,io_mem_resp_bits_rdata,io_mem_resp_bits_cmd); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_392) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec: ",_T_801); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_392) begin
          $fwrite(32'h80000002,"io.ipf:%d hitinstrPF:%d missIPF:%d pf.loadPF:%d pf.storePF:%d loadPF:%d storePF:%d\n",io_ipf,hitinstrPF,missIPF,io_pf_loadPF,io_pf_storePF,1'h0,1'h0); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module EmbeddedTLBMD(
  input          clock,
  input          reset,
  output [120:0] io_tlbmd_0,
  output [120:0] io_tlbmd_1,
  output [120:0] io_tlbmd_2,
  output [120:0] io_tlbmd_3,
  input          io_write_wen,
  input  [3:0]   io_write_waymask,
  input  [120:0] io_write_wdata,
  output         io_ready
);
`ifdef RANDOMIZE_MEM_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [120:0] tlbmd_0 [0:0]; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_0__T_data; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_0__T_addr; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_0__T_6_data; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_0__T_6_addr; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_0__T_6_mask; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_0__T_6_en; // @[EmbeddedTLB.scala 38:18]
  reg [120:0] tlbmd_1 [0:0]; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_1__T_data; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_1__T_addr; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_1__T_6_data; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_1__T_6_addr; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_1__T_6_mask; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_1__T_6_en; // @[EmbeddedTLB.scala 38:18]
  reg [120:0] tlbmd_2 [0:0]; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_2__T_data; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_2__T_addr; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_2__T_6_data; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_2__T_6_addr; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_2__T_6_mask; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_2__T_6_en; // @[EmbeddedTLB.scala 38:18]
  reg [120:0] tlbmd_3 [0:0]; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_3__T_data; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_3__T_addr; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_3__T_6_data; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_3__T_6_addr; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_3__T_6_mask; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_3__T_6_en; // @[EmbeddedTLB.scala 38:18]
  reg  resetState; // @[EmbeddedTLB.scala 42:27]
  wire  _GEN_1 = resetState ? 1'h0 : resetState; // @[EmbeddedTLB.scala 44:22]
  wire [3:0] waymask = resetState ? 4'hf : io_write_waymask; // @[EmbeddedTLB.scala 53:20]
  assign tlbmd_0__T_addr = 1'h0;
  assign tlbmd_0__T_data = tlbmd_0[tlbmd_0__T_addr]; // @[EmbeddedTLB.scala 38:18]
  assign tlbmd_0__T_6_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_0__T_6_addr = 1'h0;
  assign tlbmd_0__T_6_mask = waymask[0];
  assign tlbmd_0__T_6_en = resetState | io_write_wen;
  assign tlbmd_1__T_addr = 1'h0;
  assign tlbmd_1__T_data = tlbmd_1[tlbmd_1__T_addr]; // @[EmbeddedTLB.scala 38:18]
  assign tlbmd_1__T_6_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_1__T_6_addr = 1'h0;
  assign tlbmd_1__T_6_mask = waymask[1];
  assign tlbmd_1__T_6_en = resetState | io_write_wen;
  assign tlbmd_2__T_addr = 1'h0;
  assign tlbmd_2__T_data = tlbmd_2[tlbmd_2__T_addr]; // @[EmbeddedTLB.scala 38:18]
  assign tlbmd_2__T_6_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_2__T_6_addr = 1'h0;
  assign tlbmd_2__T_6_mask = waymask[2];
  assign tlbmd_2__T_6_en = resetState | io_write_wen;
  assign tlbmd_3__T_addr = 1'h0;
  assign tlbmd_3__T_data = tlbmd_3[tlbmd_3__T_addr]; // @[EmbeddedTLB.scala 38:18]
  assign tlbmd_3__T_6_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_3__T_6_addr = 1'h0;
  assign tlbmd_3__T_6_mask = waymask[3];
  assign tlbmd_3__T_6_en = resetState | io_write_wen;
  assign io_tlbmd_0 = tlbmd_0__T_data; // @[EmbeddedTLB.scala 39:12]
  assign io_tlbmd_1 = tlbmd_1__T_data; // @[EmbeddedTLB.scala 39:12]
  assign io_tlbmd_2 = tlbmd_2__T_data; // @[EmbeddedTLB.scala 39:12]
  assign io_tlbmd_3 = tlbmd_3__T_data; // @[EmbeddedTLB.scala 39:12]
  assign io_ready = ~resetState; // @[EmbeddedTLB.scala 59:12]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {4{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    tlbmd_0[initvar] = _RAND_0[120:0];
  _RAND_1 = {4{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    tlbmd_1[initvar] = _RAND_1[120:0];
  _RAND_2 = {4{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    tlbmd_2[initvar] = _RAND_2[120:0];
  _RAND_3 = {4{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    tlbmd_3[initvar] = _RAND_3[120:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  resetState = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(tlbmd_0__T_6_en & tlbmd_0__T_6_mask) begin
      tlbmd_0[tlbmd_0__T_6_addr] <= tlbmd_0__T_6_data; // @[EmbeddedTLB.scala 38:18]
    end
    if(tlbmd_1__T_6_en & tlbmd_1__T_6_mask) begin
      tlbmd_1[tlbmd_1__T_6_addr] <= tlbmd_1__T_6_data; // @[EmbeddedTLB.scala 38:18]
    end
    if(tlbmd_2__T_6_en & tlbmd_2__T_6_mask) begin
      tlbmd_2[tlbmd_2__T_6_addr] <= tlbmd_2__T_6_data; // @[EmbeddedTLB.scala 38:18]
    end
    if(tlbmd_3__T_6_en & tlbmd_3__T_6_mask) begin
      tlbmd_3[tlbmd_3__T_6_addr] <= tlbmd_3__T_6_data; // @[EmbeddedTLB.scala 38:18]
    end
    resetState <= reset | _GEN_1;
  end
endmodule
module EmbeddedTLB(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [38:0] io_in_req_bits_addr,
  input  [86:0] io_in_req_bits_user,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  output [86:0] io_in_resp_bits_user,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [3:0]  io_out_req_bits_cmd,
  output [63:0] io_out_req_bits_wdata,
  output [86:0] io_out_req_bits_user,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [63:0] io_out_resp_bits_rdata,
  input  [86:0] io_out_resp_bits_user,
  input         io_mem_req_ready,
  output        io_mem_req_valid,
  output [31:0] io_mem_req_bits_addr,
  output [3:0]  io_mem_req_bits_cmd,
  output [63:0] io_mem_req_bits_wdata,
  input         io_mem_resp_valid,
  input  [3:0]  io_mem_resp_bits_cmd,
  input  [63:0] io_mem_resp_bits_rdata,
  input         io_flush,
  input  [1:0]  io_csrMMU_priviledgeMode,
  output        io_csrMMU_loadPF,
  output        io_csrMMU_storePF,
  input         io_cacheEmpty,
  output        io_ipf,
  input  [63:0] CSRSATP,
  input         DISPLAY_ENABLE,
  input         MOUFlushTLB
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [95:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire  tlbExec_clock; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_reset; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_in_ready; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_in_valid; // @[EmbeddedTLB.scala 80:23]
  wire [38:0] tlbExec_io_in_bits_addr; // @[EmbeddedTLB.scala 80:23]
  wire [86:0] tlbExec_io_in_bits_user; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_out_ready; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_out_valid; // @[EmbeddedTLB.scala 80:23]
  wire [31:0] tlbExec_io_out_bits_addr; // @[EmbeddedTLB.scala 80:23]
  wire [86:0] tlbExec_io_out_bits_user; // @[EmbeddedTLB.scala 80:23]
  wire [120:0] tlbExec_io_md_0; // @[EmbeddedTLB.scala 80:23]
  wire [120:0] tlbExec_io_md_1; // @[EmbeddedTLB.scala 80:23]
  wire [120:0] tlbExec_io_md_2; // @[EmbeddedTLB.scala 80:23]
  wire [120:0] tlbExec_io_md_3; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mdWrite_wen; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mdWrite_windex; // @[EmbeddedTLB.scala 80:23]
  wire [3:0] tlbExec_io_mdWrite_waymask; // @[EmbeddedTLB.scala 80:23]
  wire [120:0] tlbExec_io_mdWrite_wdata; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mdReady; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mem_req_ready; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mem_req_valid; // @[EmbeddedTLB.scala 80:23]
  wire [31:0] tlbExec_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 80:23]
  wire [2:0] tlbExec_io_mem_req_bits_size; // @[EmbeddedTLB.scala 80:23]
  wire [3:0] tlbExec_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 80:23]
  wire [7:0] tlbExec_io_mem_req_bits_wmask; // @[EmbeddedTLB.scala 80:23]
  wire [63:0] tlbExec_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mem_resp_ready; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mem_resp_valid; // @[EmbeddedTLB.scala 80:23]
  wire [3:0] tlbExec_io_mem_resp_bits_cmd; // @[EmbeddedTLB.scala 80:23]
  wire [63:0] tlbExec_io_mem_resp_bits_rdata; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_flush; // @[EmbeddedTLB.scala 80:23]
  wire [63:0] tlbExec_io_satp; // @[EmbeddedTLB.scala 80:23]
  wire [1:0] tlbExec_io_pf_priviledgeMode; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_pf_loadPF; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_pf_storePF; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_ipf; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_isFinish; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_DISPLAY_ENABLE; // @[EmbeddedTLB.scala 80:23]
  wire  mdTLB_clock; // @[EmbeddedTLB.scala 82:21]
  wire  mdTLB_reset; // @[EmbeddedTLB.scala 82:21]
  wire [120:0] mdTLB_io_tlbmd_0; // @[EmbeddedTLB.scala 82:21]
  wire [120:0] mdTLB_io_tlbmd_1; // @[EmbeddedTLB.scala 82:21]
  wire [120:0] mdTLB_io_tlbmd_2; // @[EmbeddedTLB.scala 82:21]
  wire [120:0] mdTLB_io_tlbmd_3; // @[EmbeddedTLB.scala 82:21]
  wire  mdTLB_io_write_wen; // @[EmbeddedTLB.scala 82:21]
  wire [3:0] mdTLB_io_write_waymask; // @[EmbeddedTLB.scala 82:21]
  wire [120:0] mdTLB_io_write_wdata; // @[EmbeddedTLB.scala 82:21]
  wire  mdTLB_io_ready; // @[EmbeddedTLB.scala 82:21]
  reg [120:0] _T__0; // @[Reg.scala 15:16]
  reg [120:0] _T__1; // @[Reg.scala 15:16]
  reg [120:0] _T__2; // @[Reg.scala 15:16]
  reg [120:0] _T__3; // @[Reg.scala 15:16]
  wire  mdUpdate = io_in_req_valid & tlbExec_io_in_ready; // @[EmbeddedTLB.scala 114:26]
  wire  _T_14 = CSRSATP[63:60] == 4'h8; // @[EmbeddedTLB.scala 102:49]
  wire  _T_15 = io_csrMMU_priviledgeMode < 2'h3; // @[EmbeddedTLB.scala 102:86]
  wire  vmEnable = _T_14 & _T_15; // @[EmbeddedTLB.scala 102:57]
  reg  _T_16; // @[EmbeddedTLB.scala 105:24]
  wire  _GEN_4 = tlbExec_io_isFinish ? 1'h0 : _T_16; // @[EmbeddedTLB.scala 106:25]
  wire  _T_18 = mdUpdate & vmEnable; // @[EmbeddedTLB.scala 107:37]
  wire  _GEN_5 = _T_18 | _GEN_4; // @[EmbeddedTLB.scala 107:50]
  reg [38:0] _T_20_addr; // @[Reg.scala 15:16]
  reg [86:0] _T_20_user; // @[Reg.scala 15:16]
  wire  _T_22 = ~vmEnable; // @[EmbeddedTLB.scala 123:8]
  wire  _GEN_13 = _T_22 | io_out_req_ready; // @[EmbeddedTLB.scala 123:19]
  wire  _GEN_14 = _T_22 ? io_in_req_valid : tlbExec_io_out_valid; // @[EmbeddedTLB.scala 123:19]
  wire  _T_24 = tlbExec_io_ipf & vmEnable; // @[EmbeddedTLB.scala 152:26]
  wire  _T_25 = io_cacheEmpty & io_in_resp_ready; // @[EmbeddedTLB.scala 153:45]
  wire  _T_27 = _T_24 & io_cacheEmpty; // @[EmbeddedTLB.scala 157:38]
  reg [63:0] _T_28; // @[GTimer.scala 24:20]
  wire [63:0] _T_30 = _T_28 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_34 = ~reset; // @[Debug.scala 56:24]
  reg [63:0] _T_37; // @[GTimer.scala 24:20]
  wire [63:0] _T_39 = _T_37 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_46; // @[GTimer.scala 24:20]
  wire [63:0] _T_48 = _T_46 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_55; // @[GTimer.scala 24:20]
  wire [63:0] _T_57 = _T_55 + 64'h1; // @[GTimer.scala 25:12]
  EmbeddedTLBExec tlbExec ( // @[EmbeddedTLB.scala 80:23]
    .clock(tlbExec_clock),
    .reset(tlbExec_reset),
    .io_in_ready(tlbExec_io_in_ready),
    .io_in_valid(tlbExec_io_in_valid),
    .io_in_bits_addr(tlbExec_io_in_bits_addr),
    .io_in_bits_user(tlbExec_io_in_bits_user),
    .io_out_ready(tlbExec_io_out_ready),
    .io_out_valid(tlbExec_io_out_valid),
    .io_out_bits_addr(tlbExec_io_out_bits_addr),
    .io_out_bits_user(tlbExec_io_out_bits_user),
    .io_md_0(tlbExec_io_md_0),
    .io_md_1(tlbExec_io_md_1),
    .io_md_2(tlbExec_io_md_2),
    .io_md_3(tlbExec_io_md_3),
    .io_mdWrite_wen(tlbExec_io_mdWrite_wen),
    .io_mdWrite_windex(tlbExec_io_mdWrite_windex),
    .io_mdWrite_waymask(tlbExec_io_mdWrite_waymask),
    .io_mdWrite_wdata(tlbExec_io_mdWrite_wdata),
    .io_mdReady(tlbExec_io_mdReady),
    .io_mem_req_ready(tlbExec_io_mem_req_ready),
    .io_mem_req_valid(tlbExec_io_mem_req_valid),
    .io_mem_req_bits_addr(tlbExec_io_mem_req_bits_addr),
    .io_mem_req_bits_size(tlbExec_io_mem_req_bits_size),
    .io_mem_req_bits_cmd(tlbExec_io_mem_req_bits_cmd),
    .io_mem_req_bits_wmask(tlbExec_io_mem_req_bits_wmask),
    .io_mem_req_bits_wdata(tlbExec_io_mem_req_bits_wdata),
    .io_mem_resp_ready(tlbExec_io_mem_resp_ready),
    .io_mem_resp_valid(tlbExec_io_mem_resp_valid),
    .io_mem_resp_bits_cmd(tlbExec_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_rdata(tlbExec_io_mem_resp_bits_rdata),
    .io_flush(tlbExec_io_flush),
    .io_satp(tlbExec_io_satp),
    .io_pf_priviledgeMode(tlbExec_io_pf_priviledgeMode),
    .io_pf_loadPF(tlbExec_io_pf_loadPF),
    .io_pf_storePF(tlbExec_io_pf_storePF),
    .io_ipf(tlbExec_io_ipf),
    .io_isFinish(tlbExec_io_isFinish),
    .DISPLAY_ENABLE(tlbExec_DISPLAY_ENABLE)
  );
  EmbeddedTLBMD mdTLB ( // @[EmbeddedTLB.scala 82:21]
    .clock(mdTLB_clock),
    .reset(mdTLB_reset),
    .io_tlbmd_0(mdTLB_io_tlbmd_0),
    .io_tlbmd_1(mdTLB_io_tlbmd_1),
    .io_tlbmd_2(mdTLB_io_tlbmd_2),
    .io_tlbmd_3(mdTLB_io_tlbmd_3),
    .io_write_wen(mdTLB_io_write_wen),
    .io_write_waymask(mdTLB_io_write_waymask),
    .io_write_wdata(mdTLB_io_write_wdata),
    .io_ready(mdTLB_io_ready)
  );
  assign io_in_req_ready = _T_22 ? io_out_req_ready : tlbExec_io_in_ready; // @[EmbeddedTLB.scala 110:16 EmbeddedTLB.scala 127:21]
  assign io_in_resp_valid = _T_27 | io_out_resp_valid; // @[EmbeddedTLB.scala 138:15 EmbeddedTLB.scala 158:24]
  assign io_in_resp_bits_cmd = 4'h6; // @[EmbeddedTLB.scala 138:15 EmbeddedTLB.scala 160:27]
  assign io_in_resp_bits_rdata = _T_27 ? 64'h0 : io_out_resp_bits_rdata; // @[EmbeddedTLB.scala 138:15 EmbeddedTLB.scala 159:29]
  assign io_in_resp_bits_user = _T_27 ? tlbExec_io_in_bits_user : io_out_resp_bits_user; // @[EmbeddedTLB.scala 138:15 EmbeddedTLB.scala 161:34]
  assign io_out_req_valid = _T_24 ? 1'h0 : _GEN_14; // @[EmbeddedTLB.scala 126:22 EmbeddedTLB.scala 136:23 EmbeddedTLB.scala 154:24]
  assign io_out_req_bits_addr = _T_22 ? io_in_req_bits_addr[31:0] : tlbExec_io_out_bits_addr; // @[EmbeddedTLB.scala 128:26 EmbeddedTLB.scala 136:23]
  assign io_out_req_bits_cmd = 4'h0; // @[EmbeddedTLB.scala 130:25 EmbeddedTLB.scala 136:23]
  assign io_out_req_bits_wdata = 64'h0; // @[EmbeddedTLB.scala 132:27 EmbeddedTLB.scala 136:23]
  assign io_out_req_bits_user = _T_22 ? io_in_req_bits_user : tlbExec_io_out_bits_user; // @[EmbeddedTLB.scala 133:32 EmbeddedTLB.scala 136:23]
  assign io_out_resp_ready = io_in_resp_ready; // @[EmbeddedTLB.scala 138:15]
  assign io_mem_req_valid = tlbExec_io_mem_req_valid; // @[EmbeddedTLB.scala 87:18]
  assign io_mem_req_bits_addr = tlbExec_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 87:18]
  assign io_mem_req_bits_cmd = tlbExec_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 87:18]
  assign io_mem_req_bits_wdata = tlbExec_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 87:18]
  assign io_csrMMU_loadPF = 1'h0; // @[EmbeddedTLB.scala 88:17]
  assign io_csrMMU_storePF = 1'h0; // @[EmbeddedTLB.scala 88:17]
  assign io_ipf = _T_27 & tlbExec_io_ipf; // @[EmbeddedTLB.scala 94:10 EmbeddedTLB.scala 162:14]
  assign tlbExec_clock = clock;
  assign tlbExec_reset = reset;
  assign tlbExec_io_in_valid = _T_16; // @[EmbeddedTLB.scala 112:17]
  assign tlbExec_io_in_bits_addr = _T_20_addr; // @[EmbeddedTLB.scala 111:16]
  assign tlbExec_io_in_bits_user = _T_20_user; // @[EmbeddedTLB.scala 111:16]
  assign tlbExec_io_out_ready = _T_24 ? _T_25 : _GEN_13; // @[EmbeddedTLB.scala 124:26 EmbeddedTLB.scala 136:23 EmbeddedTLB.scala 153:28]
  assign tlbExec_io_md_0 = _T__0; // @[EmbeddedTLB.scala 89:17]
  assign tlbExec_io_md_1 = _T__1; // @[EmbeddedTLB.scala 89:17]
  assign tlbExec_io_md_2 = _T__2; // @[EmbeddedTLB.scala 89:17]
  assign tlbExec_io_md_3 = _T__3; // @[EmbeddedTLB.scala 89:17]
  assign tlbExec_io_mdReady = mdTLB_io_ready; // @[EmbeddedTLB.scala 90:22]
  assign tlbExec_io_mem_req_ready = io_mem_req_ready; // @[EmbeddedTLB.scala 87:18]
  assign tlbExec_io_mem_resp_valid = io_mem_resp_valid; // @[EmbeddedTLB.scala 87:18]
  assign tlbExec_io_mem_resp_bits_cmd = io_mem_resp_bits_cmd; // @[EmbeddedTLB.scala 87:18]
  assign tlbExec_io_mem_resp_bits_rdata = io_mem_resp_bits_rdata; // @[EmbeddedTLB.scala 87:18]
  assign tlbExec_io_flush = io_flush; // @[EmbeddedTLB.scala 85:20]
  assign tlbExec_io_satp = CSRSATP; // @[EmbeddedTLB.scala 86:19]
  assign tlbExec_io_pf_priviledgeMode = io_csrMMU_priviledgeMode; // @[EmbeddedTLB.scala 88:17]
  assign tlbExec_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign mdTLB_clock = clock;
  assign mdTLB_reset = reset | MOUFlushTLB; // @[EmbeddedTLB.scala 99:15]
  assign mdTLB_io_write_wen = tlbExec_io_mdWrite_wen; // @[EmbeddedTLB.scala 92:18]
  assign mdTLB_io_write_waymask = tlbExec_io_mdWrite_waymask; // @[EmbeddedTLB.scala 92:18]
  assign mdTLB_io_write_wdata = tlbExec_io_mdWrite_wdata; // @[EmbeddedTLB.scala 92:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  _T__0 = _RAND_0[120:0];
  _RAND_1 = {4{`RANDOM}};
  _T__1 = _RAND_1[120:0];
  _RAND_2 = {4{`RANDOM}};
  _T__2 = _RAND_2[120:0];
  _RAND_3 = {4{`RANDOM}};
  _T__3 = _RAND_3[120:0];
  _RAND_4 = {1{`RANDOM}};
  _T_16 = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  _T_20_addr = _RAND_5[38:0];
  _RAND_6 = {3{`RANDOM}};
  _T_20_user = _RAND_6[86:0];
  _RAND_7 = {2{`RANDOM}};
  _T_28 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  _T_37 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  _T_46 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  _T_55 = _RAND_10[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (mdUpdate) begin
      _T__0 <= mdTLB_io_tlbmd_0;
    end
    if (mdUpdate) begin
      _T__1 <= mdTLB_io_tlbmd_1;
    end
    if (mdUpdate) begin
      _T__2 <= mdTLB_io_tlbmd_2;
    end
    if (mdUpdate) begin
      _T__3 <= mdTLB_io_tlbmd_3;
    end
    if (reset) begin
      _T_16 <= 1'h0;
    end else if (io_flush) begin
      _T_16 <= 1'h0;
    end else begin
      _T_16 <= _GEN_5;
    end
    if (mdUpdate) begin
      _T_20_addr <= io_in_req_bits_addr;
    end
    if (mdUpdate) begin
      _T_20_user <= io_in_req_bits_user;
    end
    if (reset) begin
      _T_28 <= 64'h0;
    end else begin
      _T_28 <= _T_30;
    end
    if (reset) begin
      _T_37 <= 64'h0;
    end else begin
      _T_37 <= _T_39;
    end
    if (reset) begin
      _T_46 <= 64'h0;
    end else begin
      _T_46 <= _T_48;
    end
    if (reset) begin
      _T_55 <= 64'h0;
    end else begin
      _T_55 <= _T_57;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_34) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLB: ",_T_28); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_34) begin
          $fwrite(32'h80000002,"InReq(%d, %d) InResp(%d, %d) OutReq(%d, %d) OutResp(%d, %d) vmEnable:%d mode:%d\n",io_in_req_valid,io_in_req_ready,io_in_resp_valid,io_in_resp_ready,io_out_req_valid,io_out_req_ready,io_out_resp_valid,io_out_resp_ready,vmEnable,io_csrMMU_priviledgeMode); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_34) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLB: ",_T_37); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_34) begin
          $fwrite(32'h80000002,"InReq: addr:%x cmd:%d wdata:%x OutReq: addr:%x cmd:%x wdata:%x\n",io_in_req_bits_addr,4'h0,64'h0,io_out_req_bits_addr,io_out_req_bits_cmd,io_out_req_bits_wdata); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_34) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLB: ",_T_46); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_34) begin
          $fwrite(32'h80000002,"OutResp: rdata:%x cmd:%x Inresp: rdata:%x cmd:%x\n",io_out_resp_bits_rdata,4'h6,io_in_resp_bits_rdata,io_in_resp_bits_cmd); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_34) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLB: ",_T_55); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_34) begin
          $fwrite(32'h80000002,"satp:%x flush:%d cacheEmpty:%d instrPF:%d loadPF:%d storePF:%d \n",CSRSATP,io_flush,io_cacheEmpty,io_ipf,io_csrMMU_loadPF,io_csrMMU_storePF); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CacheStage1(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [2:0]  io_in_bits_size,
  input  [3:0]  io_in_bits_cmd,
  input  [7:0]  io_in_bits_wmask,
  input  [63:0] io_in_bits_wdata,
  input  [86:0] io_in_bits_user,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_req_addr,
  output [86:0] io_out_bits_req_user,
  input         io_metaReadBus_req_ready,
  output        io_metaReadBus_req_valid,
  output [6:0]  io_metaReadBus_req_bits_setIdx,
  input  [18:0] io_metaReadBus_resp_data_0_tag,
  input         io_metaReadBus_resp_data_0_valid,
  input         io_metaReadBus_resp_data_0_dirty,
  input  [18:0] io_metaReadBus_resp_data_1_tag,
  input         io_metaReadBus_resp_data_1_valid,
  input         io_metaReadBus_resp_data_1_dirty,
  input  [18:0] io_metaReadBus_resp_data_2_tag,
  input         io_metaReadBus_resp_data_2_valid,
  input         io_metaReadBus_resp_data_2_dirty,
  input  [18:0] io_metaReadBus_resp_data_3_tag,
  input         io_metaReadBus_resp_data_3_valid,
  input         io_metaReadBus_resp_data_3_dirty,
  input         io_dataReadBus_req_ready,
  output        io_dataReadBus_req_valid,
  output [9:0]  io_dataReadBus_req_bits_setIdx,
  input  [63:0] io_dataReadBus_resp_data_0_data,
  input  [63:0] io_dataReadBus_resp_data_1_data,
  input  [63:0] io_dataReadBus_resp_data_2_data,
  input  [63:0] io_dataReadBus_resp_data_3_data,
  input         DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  _T = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  reg [63:0] _T_7; // @[GTimer.scala 24:20]
  wire [63:0] _T_9 = _T_7 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_11 = _T & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  wire  _T_13 = ~reset; // @[Debug.scala 56:24]
  wire  _T_35 = io_in_valid & io_metaReadBus_req_ready; // @[Cache.scala 133:31]
  wire  _T_37 = ~io_in_valid; // @[Cache.scala 134:19]
  wire  _T_38 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_39 = _T_37 | _T_38; // @[Cache.scala 134:32]
  wire  _T_40 = _T_39 & io_metaReadBus_req_ready; // @[Cache.scala 134:50]
  reg [63:0] _T_42; // @[GTimer.scala 24:20]
  wire [63:0] _T_44 = _T_42 + 64'h1; // @[GTimer.scala 25:12]
  assign io_in_ready = _T_40 & io_dataReadBus_req_ready; // @[Cache.scala 134:15]
  assign io_out_valid = _T_35 & io_dataReadBus_req_ready; // @[Cache.scala 133:16]
  assign io_out_bits_req_addr = io_in_bits_addr; // @[Cache.scala 132:19]
  assign io_out_bits_req_user = io_in_bits_user; // @[Cache.scala 132:19]
  assign io_metaReadBus_req_valid = io_in_valid & io_out_ready; // @[SRAMTemplate.scala 53:20]
  assign io_metaReadBus_req_bits_setIdx = io_in_bits_addr[12:6]; // @[SRAMTemplate.scala 26:17]
  assign io_dataReadBus_req_valid = io_in_valid & io_out_ready; // @[SRAMTemplate.scala 53:20]
  assign io_dataReadBus_req_bits_setIdx = {io_in_bits_addr[12:6],io_in_bits_addr[5:3]}; // @[SRAMTemplate.scala 26:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  _T_7 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  _T_42 = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_7 <= 64'h0;
    end else begin
      _T_7 <= _T_9;
    end
    if (reset) begin
      _T_42 <= 64'h0;
    end else begin
      _T_42 <= _T_44;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_11 & _T_13) begin
          $fwrite(32'h80000002,"[%d] CacheStage1: ",_T_7); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_11 & _T_13) begin
          $fwrite(32'h80000002,"[L1$] cache stage1, addr in: %x, user: %x id: %x\n",io_in_bits_addr,io_in_bits_user,1'h0); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_13) begin
          $fwrite(32'h80000002,"[%d] CacheStage1: ",_T_42); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_13) begin
          $fwrite(32'h80000002,"in.ready = %d, in.valid = %d, out.valid = %d, out.ready = %d, addr = %x, cmd = %x, dataReadBus.req.valid = %d\n",io_in_ready,io_in_valid,io_out_valid,io_out_ready,io_in_bits_addr,4'h0,io_dataReadBus_req_valid); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CacheStage2(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_req_addr,
  input  [2:0]  io_in_bits_req_size,
  input  [3:0]  io_in_bits_req_cmd,
  input  [7:0]  io_in_bits_req_wmask,
  input  [63:0] io_in_bits_req_wdata,
  input  [86:0] io_in_bits_req_user,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_req_addr,
  output [86:0] io_out_bits_req_user,
  output [18:0] io_out_bits_metas_0_tag,
  output        io_out_bits_metas_0_valid,
  output        io_out_bits_metas_0_dirty,
  output [18:0] io_out_bits_metas_1_tag,
  output        io_out_bits_metas_1_valid,
  output        io_out_bits_metas_1_dirty,
  output [18:0] io_out_bits_metas_2_tag,
  output        io_out_bits_metas_2_valid,
  output        io_out_bits_metas_2_dirty,
  output [18:0] io_out_bits_metas_3_tag,
  output        io_out_bits_metas_3_valid,
  output        io_out_bits_metas_3_dirty,
  output [63:0] io_out_bits_datas_0_data,
  output [63:0] io_out_bits_datas_1_data,
  output [63:0] io_out_bits_datas_2_data,
  output [63:0] io_out_bits_datas_3_data,
  output        io_out_bits_hit,
  output [3:0]  io_out_bits_waymask,
  output        io_out_bits_mmio,
  output        io_out_bits_isForwardData,
  output [63:0] io_out_bits_forwardData_data_data,
  output [3:0]  io_out_bits_forwardData_waymask,
  input  [18:0] io_metaReadResp_0_tag,
  input         io_metaReadResp_0_valid,
  input         io_metaReadResp_0_dirty,
  input  [18:0] io_metaReadResp_1_tag,
  input         io_metaReadResp_1_valid,
  input         io_metaReadResp_1_dirty,
  input  [18:0] io_metaReadResp_2_tag,
  input         io_metaReadResp_2_valid,
  input         io_metaReadResp_2_dirty,
  input  [18:0] io_metaReadResp_3_tag,
  input         io_metaReadResp_3_valid,
  input         io_metaReadResp_3_dirty,
  input  [63:0] io_dataReadResp_0_data,
  input  [63:0] io_dataReadResp_1_data,
  input  [63:0] io_dataReadResp_2_data,
  input  [63:0] io_dataReadResp_3_data,
  input         io_metaWriteBus_req_valid,
  input  [6:0]  io_metaWriteBus_req_bits_setIdx,
  input  [18:0] io_metaWriteBus_req_bits_data_tag,
  input         io_metaWriteBus_req_bits_data_dirty,
  input  [3:0]  io_metaWriteBus_req_bits_waymask,
  input         io_dataWriteBus_req_valid,
  input  [9:0]  io_dataWriteBus_req_bits_setIdx,
  input  [63:0] io_dataWriteBus_req_bits_data_data,
  input  [3:0]  io_dataWriteBus_req_bits_waymask,
  input         DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[Cache.scala 162:31]
  wire [6:0] addr_index = io_in_bits_req_addr[12:6]; // @[Cache.scala 162:31]
  wire [18:0] addr_tag = io_in_bits_req_addr[31:13]; // @[Cache.scala 162:31]
  wire  _T_5 = io_in_valid & io_metaWriteBus_req_valid; // @[Cache.scala 164:35]
  wire  _T_12 = io_metaWriteBus_req_bits_setIdx == addr_index; // @[Cache.scala 164:99]
  wire  isForwardMeta = _T_5 & _T_12; // @[Cache.scala 164:64]
  reg  isForwardMetaReg; // @[Cache.scala 165:33]
  wire  _GEN_0 = isForwardMeta | isForwardMetaReg; // @[Cache.scala 166:24]
  wire  _T_13 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire  _T_14 = ~io_in_valid; // @[Cache.scala 167:25]
  wire  _T_15 = _T_13 | _T_14; // @[Cache.scala 167:22]
  reg [18:0] forwardMetaReg_data_tag; // @[Reg.scala 15:16]
  reg  forwardMetaReg_data_dirty; // @[Reg.scala 15:16]
  reg [3:0] forwardMetaReg_waymask; // @[Reg.scala 15:16]
  wire [3:0] _GEN_2 = isForwardMeta ? io_metaWriteBus_req_bits_waymask : forwardMetaReg_waymask; // @[Reg.scala 16:19]
  wire  _GEN_3 = isForwardMeta ? io_metaWriteBus_req_bits_data_dirty : forwardMetaReg_data_dirty; // @[Reg.scala 16:19]
  wire [18:0] _GEN_5 = isForwardMeta ? io_metaWriteBus_req_bits_data_tag : forwardMetaReg_data_tag; // @[Reg.scala 16:19]
  wire  pickForwardMeta = isForwardMetaReg | isForwardMeta; // @[Cache.scala 171:42]
  wire  forwardWaymask_0 = _GEN_2[0]; // @[Cache.scala 173:61]
  wire  forwardWaymask_1 = _GEN_2[1]; // @[Cache.scala 173:61]
  wire  forwardWaymask_2 = _GEN_2[2]; // @[Cache.scala 173:61]
  wire  forwardWaymask_3 = _GEN_2[3]; // @[Cache.scala 173:61]
  wire  _T_16 = pickForwardMeta & forwardWaymask_0; // @[Cache.scala 175:39]
  wire [18:0] metaWay_0_tag = _T_16 ? _GEN_5 : io_metaReadResp_0_tag; // @[Cache.scala 175:22]
  wire  metaWay_0_valid = _T_16 | io_metaReadResp_0_valid; // @[Cache.scala 175:22]
  wire  _T_18 = pickForwardMeta & forwardWaymask_1; // @[Cache.scala 175:39]
  wire [18:0] metaWay_1_tag = _T_18 ? _GEN_5 : io_metaReadResp_1_tag; // @[Cache.scala 175:22]
  wire  metaWay_1_valid = _T_18 | io_metaReadResp_1_valid; // @[Cache.scala 175:22]
  wire  _T_20 = pickForwardMeta & forwardWaymask_2; // @[Cache.scala 175:39]
  wire [18:0] metaWay_2_tag = _T_20 ? _GEN_5 : io_metaReadResp_2_tag; // @[Cache.scala 175:22]
  wire  metaWay_2_valid = _T_20 | io_metaReadResp_2_valid; // @[Cache.scala 175:22]
  wire  _T_22 = pickForwardMeta & forwardWaymask_3; // @[Cache.scala 175:39]
  wire [18:0] metaWay_3_tag = _T_22 ? _GEN_5 : io_metaReadResp_3_tag; // @[Cache.scala 175:22]
  wire  metaWay_3_valid = _T_22 | io_metaReadResp_3_valid; // @[Cache.scala 175:22]
  wire  _T_24 = metaWay_0_tag == addr_tag; // @[Cache.scala 178:59]
  wire  _T_25 = metaWay_0_valid & _T_24; // @[Cache.scala 178:49]
  wire  _T_26 = _T_25 & io_in_valid; // @[Cache.scala 178:73]
  wire  _T_27 = metaWay_1_tag == addr_tag; // @[Cache.scala 178:59]
  wire  _T_28 = metaWay_1_valid & _T_27; // @[Cache.scala 178:49]
  wire  _T_29 = _T_28 & io_in_valid; // @[Cache.scala 178:73]
  wire  _T_30 = metaWay_2_tag == addr_tag; // @[Cache.scala 178:59]
  wire  _T_31 = metaWay_2_valid & _T_30; // @[Cache.scala 178:49]
  wire  _T_32 = _T_31 & io_in_valid; // @[Cache.scala 178:73]
  wire  _T_33 = metaWay_3_tag == addr_tag; // @[Cache.scala 178:59]
  wire  _T_34 = metaWay_3_valid & _T_33; // @[Cache.scala 178:49]
  wire  _T_35 = _T_34 & io_in_valid; // @[Cache.scala 178:73]
  wire [3:0] hitVec = {_T_35,_T_32,_T_29,_T_26}; // @[Cache.scala 178:90]
  reg [63:0] _T_39; // @[LFSR64.scala 25:23]
  wire  _T_42 = _T_39[0] ^ _T_39[1]; // @[LFSR64.scala 26:23]
  wire  _T_44 = _T_42 ^ _T_39[3]; // @[LFSR64.scala 26:33]
  wire  _T_46 = _T_44 ^ _T_39[4]; // @[LFSR64.scala 26:43]
  wire  _T_47 = _T_39 == 64'h0; // @[LFSR64.scala 28:24]
  wire [63:0] _T_49 = {_T_46,_T_39[63:1]}; // @[Cat.scala 29:58]
  wire [3:0] victimWaymask = 4'h1 << _T_39[1:0]; // @[Cache.scala 179:42]
  wire  _T_52 = ~metaWay_0_valid; // @[Cache.scala 181:45]
  wire  _T_53 = ~metaWay_1_valid; // @[Cache.scala 181:45]
  wire  _T_54 = ~metaWay_2_valid; // @[Cache.scala 181:45]
  wire  _T_55 = ~metaWay_3_valid; // @[Cache.scala 181:45]
  wire [3:0] invalidVec = {_T_55,_T_54,_T_53,_T_52}; // @[Cache.scala 181:56]
  wire  hasInvalidWay = |invalidVec; // @[Cache.scala 182:34]
  wire  _T_59 = invalidVec >= 4'h8; // @[Cache.scala 183:45]
  wire  _T_60 = invalidVec >= 4'h4; // @[Cache.scala 184:20]
  wire  _T_61 = invalidVec >= 4'h2; // @[Cache.scala 185:20]
  wire [1:0] _T_62 = _T_61 ? 2'h2 : 2'h1; // @[Cache.scala 185:8]
  wire [2:0] _T_63 = _T_60 ? 3'h4 : {{1'd0}, _T_62}; // @[Cache.scala 184:8]
  wire [3:0] refillInvalidWaymask = _T_59 ? 4'h8 : {{1'd0}, _T_63}; // @[Cache.scala 183:33]
  wire [3:0] _T_64 = hasInvalidWay ? refillInvalidWaymask : victimWaymask; // @[Cache.scala 188:49]
  wire [3:0] waymask = io_out_bits_hit ? hitVec : _T_64; // @[Cache.scala 188:20]
  wire [1:0] _T_69 = waymask[0] + waymask[1]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_71 = waymask[2] + waymask[3]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_73 = _T_69 + _T_71; // @[Bitwise.scala 47:55]
  wire  _T_75 = _T_73 > 3'h1; // @[Cache.scala 189:26]
  reg [63:0] _T_76; // @[GTimer.scala 24:20]
  wire [63:0] _T_78 = _T_76 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_82 = ~reset; // @[Debug.scala 56:24]
  reg [63:0] _T_85; // @[GTimer.scala 24:20]
  wire [63:0] _T_87 = _T_85 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_94; // @[GTimer.scala 24:20]
  wire [63:0] _T_96 = _T_94 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_103; // @[GTimer.scala 24:20]
  wire [63:0] _T_105 = _T_103 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_112; // @[GTimer.scala 24:20]
  wire [63:0] _T_114 = _T_112 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_121; // @[GTimer.scala 24:20]
  wire [63:0] _T_123 = _T_121 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_130; // @[GTimer.scala 24:20]
  wire [63:0] _T_132 = _T_130 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_139; // @[GTimer.scala 24:20]
  wire [63:0] _T_141 = _T_139 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_148; // @[GTimer.scala 24:20]
  wire [63:0] _T_150 = _T_148 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_157; // @[GTimer.scala 24:20]
  wire [63:0] _T_159 = _T_157 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_177; // @[GTimer.scala 24:20]
  wire [63:0] _T_179 = _T_177 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_197 = io_in_valid & _T_75; // @[Cache.scala 196:24]
  wire  _T_198 = ~_T_197; // @[Cache.scala 196:10]
  wire  _T_200 = _T_198 | reset; // @[Cache.scala 196:9]
  wire  _T_201 = ~_T_200; // @[Cache.scala 196:9]
  wire  _T_202 = |hitVec; // @[Cache.scala 199:44]
  wire [31:0] _T_204 = io_in_bits_req_addr ^ 32'h30000000; // @[NutCore.scala 86:11]
  wire  _T_206 = _T_204[31:28] == 4'h0; // @[NutCore.scala 86:44]
  wire [31:0] _T_207 = io_in_bits_req_addr ^ 32'h40000000; // @[NutCore.scala 86:11]
  wire  _T_209 = _T_207[31:30] == 2'h0; // @[NutCore.scala 86:44]
  wire [9:0] _T_223 = {addr_index,addr_wordIndex}; // @[Cat.scala 29:58]
  wire  _T_224 = io_dataWriteBus_req_bits_setIdx == _T_223; // @[Cache.scala 205:30]
  wire  _T_225 = io_dataWriteBus_req_valid & _T_224; // @[Cache.scala 205:13]
  wire  isForwardData = io_in_valid & _T_225; // @[Cache.scala 204:35]
  reg  isForwardDataReg; // @[Cache.scala 207:33]
  wire  _GEN_8 = isForwardData | isForwardDataReg; // @[Cache.scala 208:24]
  reg [63:0] forwardDataReg_data_data; // @[Reg.scala 15:16]
  reg [3:0] forwardDataReg_waymask; // @[Reg.scala 15:16]
  wire  _T_232 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  reg [63:0] _T_235; // @[GTimer.scala 24:20]
  wire [63:0] _T_237 = _T_235 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_250; // @[GTimer.scala 24:20]
  wire [63:0] _T_252 = _T_250 + 64'h1; // @[GTimer.scala 25:12]
  wire  _GEN_13 = _T_75 & DISPLAY_ENABLE; // @[Debug.scala 56:24]
  assign io_in_ready = _T_14 | _T_232; // @[Cache.scala 216:15]
  assign io_out_valid = io_in_valid; // @[Cache.scala 215:16]
  assign io_out_bits_req_addr = io_in_bits_req_addr; // @[Cache.scala 214:19]
  assign io_out_bits_req_user = io_in_bits_req_user; // @[Cache.scala 214:19]
  assign io_out_bits_metas_0_tag = _T_16 ? _GEN_5 : io_metaReadResp_0_tag; // @[Cache.scala 198:21]
  assign io_out_bits_metas_0_valid = _T_16 | io_metaReadResp_0_valid; // @[Cache.scala 198:21]
  assign io_out_bits_metas_0_dirty = _T_16 ? _GEN_3 : io_metaReadResp_0_dirty; // @[Cache.scala 198:21]
  assign io_out_bits_metas_1_tag = _T_18 ? _GEN_5 : io_metaReadResp_1_tag; // @[Cache.scala 198:21]
  assign io_out_bits_metas_1_valid = _T_18 | io_metaReadResp_1_valid; // @[Cache.scala 198:21]
  assign io_out_bits_metas_1_dirty = _T_18 ? _GEN_3 : io_metaReadResp_1_dirty; // @[Cache.scala 198:21]
  assign io_out_bits_metas_2_tag = _T_20 ? _GEN_5 : io_metaReadResp_2_tag; // @[Cache.scala 198:21]
  assign io_out_bits_metas_2_valid = _T_20 | io_metaReadResp_2_valid; // @[Cache.scala 198:21]
  assign io_out_bits_metas_2_dirty = _T_20 ? _GEN_3 : io_metaReadResp_2_dirty; // @[Cache.scala 198:21]
  assign io_out_bits_metas_3_tag = _T_22 ? _GEN_5 : io_metaReadResp_3_tag; // @[Cache.scala 198:21]
  assign io_out_bits_metas_3_valid = _T_22 | io_metaReadResp_3_valid; // @[Cache.scala 198:21]
  assign io_out_bits_metas_3_dirty = _T_22 ? _GEN_3 : io_metaReadResp_3_dirty; // @[Cache.scala 198:21]
  assign io_out_bits_datas_0_data = io_dataReadResp_0_data; // @[Cache.scala 201:21]
  assign io_out_bits_datas_1_data = io_dataReadResp_1_data; // @[Cache.scala 201:21]
  assign io_out_bits_datas_2_data = io_dataReadResp_2_data; // @[Cache.scala 201:21]
  assign io_out_bits_datas_3_data = io_dataReadResp_3_data; // @[Cache.scala 201:21]
  assign io_out_bits_hit = io_in_valid & _T_202; // @[Cache.scala 199:19]
  assign io_out_bits_waymask = io_out_bits_hit ? hitVec : _T_64; // @[Cache.scala 200:23]
  assign io_out_bits_mmio = _T_206 | _T_209; // @[Cache.scala 202:20]
  assign io_out_bits_isForwardData = isForwardDataReg | isForwardData; // @[Cache.scala 211:29]
  assign io_out_bits_forwardData_data_data = isForwardData ? io_dataWriteBus_req_bits_data_data : forwardDataReg_data_data; // @[Cache.scala 212:27]
  assign io_out_bits_forwardData_waymask = isForwardData ? io_dataWriteBus_req_bits_waymask : forwardDataReg_waymask; // @[Cache.scala 212:27]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  isForwardMetaReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  forwardMetaReg_data_tag = _RAND_1[18:0];
  _RAND_2 = {1{`RANDOM}};
  forwardMetaReg_data_dirty = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  forwardMetaReg_waymask = _RAND_3[3:0];
  _RAND_4 = {2{`RANDOM}};
  _T_39 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  _T_76 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  _T_85 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  _T_94 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  _T_103 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  _T_112 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  _T_121 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  _T_130 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  _T_139 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  _T_148 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  _T_157 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  _T_177 = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  isForwardDataReg = _RAND_16[0:0];
  _RAND_17 = {2{`RANDOM}};
  forwardDataReg_data_data = _RAND_17[63:0];
  _RAND_18 = {1{`RANDOM}};
  forwardDataReg_waymask = _RAND_18[3:0];
  _RAND_19 = {2{`RANDOM}};
  _T_235 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  _T_250 = _RAND_20[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      isForwardMetaReg <= 1'h0;
    end else if (_T_15) begin
      isForwardMetaReg <= 1'h0;
    end else begin
      isForwardMetaReg <= _GEN_0;
    end
    if (isForwardMeta) begin
      forwardMetaReg_data_tag <= io_metaWriteBus_req_bits_data_tag;
    end
    if (isForwardMeta) begin
      forwardMetaReg_data_dirty <= io_metaWriteBus_req_bits_data_dirty;
    end
    if (isForwardMeta) begin
      forwardMetaReg_waymask <= io_metaWriteBus_req_bits_waymask;
    end
    if (reset) begin
      _T_39 <= 64'h1234567887654321;
    end else if (_T_47) begin
      _T_39 <= 64'h1;
    end else begin
      _T_39 <= _T_49;
    end
    if (reset) begin
      _T_76 <= 64'h0;
    end else begin
      _T_76 <= _T_78;
    end
    if (reset) begin
      _T_85 <= 64'h0;
    end else begin
      _T_85 <= _T_87;
    end
    if (reset) begin
      _T_94 <= 64'h0;
    end else begin
      _T_94 <= _T_96;
    end
    if (reset) begin
      _T_103 <= 64'h0;
    end else begin
      _T_103 <= _T_105;
    end
    if (reset) begin
      _T_112 <= 64'h0;
    end else begin
      _T_112 <= _T_114;
    end
    if (reset) begin
      _T_121 <= 64'h0;
    end else begin
      _T_121 <= _T_123;
    end
    if (reset) begin
      _T_130 <= 64'h0;
    end else begin
      _T_130 <= _T_132;
    end
    if (reset) begin
      _T_139 <= 64'h0;
    end else begin
      _T_139 <= _T_141;
    end
    if (reset) begin
      _T_148 <= 64'h0;
    end else begin
      _T_148 <= _T_150;
    end
    if (reset) begin
      _T_157 <= 64'h0;
    end else begin
      _T_157 <= _T_159;
    end
    if (reset) begin
      _T_177 <= 64'h0;
    end else begin
      _T_177 <= _T_179;
    end
    if (reset) begin
      isForwardDataReg <= 1'h0;
    end else if (_T_15) begin
      isForwardDataReg <= 1'h0;
    end else begin
      isForwardDataReg <= _GEN_8;
    end
    if (isForwardData) begin
      forwardDataReg_data_data <= io_dataWriteBus_req_bits_data_data;
    end
    if (isForwardData) begin
      forwardDataReg_waymask <= io_dataWriteBus_req_bits_waymask;
    end
    if (reset) begin
      _T_235 <= 64'h0;
    end else begin
      _T_235 <= _T_237;
    end
    if (reset) begin
      _T_250 <= 64'h0;
    end else begin
      _T_250 <= _T_252;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2: ",_T_76); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] metaWay %x metat %x reqt %x\n",metaWay_0_valid,metaWay_0_tag,addr_tag); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2: ",_T_85); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] metaWay %x metat %x reqt %x\n",metaWay_1_valid,metaWay_1_tag,addr_tag); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2: ",_T_94); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] metaWay %x metat %x reqt %x\n",metaWay_2_valid,metaWay_2_tag,addr_tag); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2: ",_T_103); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] metaWay %x metat %x reqt %x\n",metaWay_3_valid,metaWay_3_tag,addr_tag); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2: ",_T_112); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] metaReadResp %x metat %x reqt %x\n",io_metaReadResp_0_valid,io_metaReadResp_0_tag,addr_tag); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2: ",_T_121); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] metaReadResp %x metat %x reqt %x\n",io_metaReadResp_1_valid,io_metaReadResp_1_tag,addr_tag); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2: ",_T_130); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] metaReadResp %x metat %x reqt %x\n",io_metaReadResp_2_valid,io_metaReadResp_2_tag,addr_tag); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2: ",_T_139); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] metaReadResp %x metat %x reqt %x\n",io_metaReadResp_3_valid,io_metaReadResp_3_tag,addr_tag); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2: ",_T_148); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] forwardMetaReg isForwardMetaReg %x %x metat %x wm %b\n",isForwardMetaReg,1'h1,forwardMetaReg_data_tag,forwardMetaReg_waymask); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2: ",_T_157); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] forwardMeta isForwardMeta %x %x metat %x wm %b\n",isForwardMeta,1'h1,io_metaWriteBus_req_bits_data_tag,io_metaWriteBus_req_bits_waymask); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2: ",_T_177); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] hit %b wmask %b hitvec %b\n",io_out_bits_hit,_GEN_2,hitVec); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_201) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Cache.scala:196 assert(!(io.in.valid && PopCount(waymask) > 1.U))\n"); // @[Cache.scala 196:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_201) begin
          $fatal; // @[Cache.scala 196:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2: ",_T_235); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_82) begin
          $fwrite(32'h80000002,"[isFD:%d isFDreg:%d inFire:%d invalid:%d \n",isForwardData,isForwardDataReg,_T_13,io_in_valid); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2: ",_T_250); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_82) begin
          $fwrite(32'h80000002,"[isFM:%d isFMreg:%d metawreq:%x widx:%x ridx:%x \n",isForwardMeta,isForwardMetaReg,io_metaWriteBus_req_valid,io_metaWriteBus_req_bits_setIdx,addr_index); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Arbiter(
  input         io_in_0_valid,
  input  [6:0]  io_in_0_bits_setIdx,
  input  [18:0] io_in_0_bits_data_tag,
  input         io_in_0_bits_data_dirty,
  input  [3:0]  io_in_0_bits_waymask,
  input         io_in_1_valid,
  input  [6:0]  io_in_1_bits_setIdx,
  input  [18:0] io_in_1_bits_data_tag,
  input         io_in_1_bits_data_dirty,
  input  [3:0]  io_in_1_bits_waymask,
  output        io_out_valid,
  output [6:0]  io_out_bits_setIdx,
  output [18:0] io_out_bits_data_tag,
  output        io_out_bits_data_dirty,
  output [3:0]  io_out_bits_waymask
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  wire  _T_2 = ~grant_1; // @[Arbiter.scala 135:19]
  assign io_out_valid = _T_2 | io_in_1_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_data_tag = io_in_0_valid ? io_in_0_bits_data_tag : io_in_1_bits_data_tag; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_data_dirty = io_in_0_valid ? io_in_0_bits_data_dirty : io_in_1_bits_data_dirty; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_waymask = io_in_0_valid ? io_in_0_bits_waymask : io_in_1_bits_waymask; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
endmodule
module Arbiter_1(
  input         io_in_0_valid,
  input  [9:0]  io_in_0_bits_setIdx,
  input  [63:0] io_in_0_bits_data_data,
  input  [3:0]  io_in_0_bits_waymask,
  input         io_in_1_valid,
  input  [9:0]  io_in_1_bits_setIdx,
  input  [63:0] io_in_1_bits_data_data,
  input  [3:0]  io_in_1_bits_waymask,
  output        io_out_valid,
  output [9:0]  io_out_bits_setIdx,
  output [63:0] io_out_bits_data_data,
  output [3:0]  io_out_bits_waymask
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  wire  _T_2 = ~grant_1; // @[Arbiter.scala 135:19]
  assign io_out_valid = _T_2 | io_in_1_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_data_data = io_in_0_valid ? io_in_0_bits_data_data : io_in_1_bits_data_data; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_waymask = io_in_0_valid ? io_in_0_bits_waymask : io_in_1_bits_waymask; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
endmodule
module CacheStage3(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_req_addr,
  input  [2:0]  io_in_bits_req_size,
  input  [3:0]  io_in_bits_req_cmd,
  input  [7:0]  io_in_bits_req_wmask,
  input  [63:0] io_in_bits_req_wdata,
  input  [86:0] io_in_bits_req_user,
  input  [18:0] io_in_bits_metas_0_tag,
  input         io_in_bits_metas_0_valid,
  input         io_in_bits_metas_0_dirty,
  input  [18:0] io_in_bits_metas_1_tag,
  input         io_in_bits_metas_1_valid,
  input         io_in_bits_metas_1_dirty,
  input  [18:0] io_in_bits_metas_2_tag,
  input         io_in_bits_metas_2_valid,
  input         io_in_bits_metas_2_dirty,
  input  [18:0] io_in_bits_metas_3_tag,
  input         io_in_bits_metas_3_valid,
  input         io_in_bits_metas_3_dirty,
  input  [63:0] io_in_bits_datas_0_data,
  input  [63:0] io_in_bits_datas_1_data,
  input  [63:0] io_in_bits_datas_2_data,
  input  [63:0] io_in_bits_datas_3_data,
  input         io_in_bits_hit,
  input  [3:0]  io_in_bits_waymask,
  input         io_in_bits_mmio,
  input         io_in_bits_isForwardData,
  input  [63:0] io_in_bits_forwardData_data_data,
  input  [3:0]  io_in_bits_forwardData_waymask,
  input         io_out_ready,
  output        io_out_valid,
  output [3:0]  io_out_bits_cmd,
  output [63:0] io_out_bits_rdata,
  output [86:0] io_out_bits_user,
  output        io_isFinish,
  input         io_flush,
  input         io_dataReadBus_req_ready,
  output        io_dataReadBus_req_valid,
  output [9:0]  io_dataReadBus_req_bits_setIdx,
  input  [63:0] io_dataReadBus_resp_data_0_data,
  input  [63:0] io_dataReadBus_resp_data_1_data,
  input  [63:0] io_dataReadBus_resp_data_2_data,
  input  [63:0] io_dataReadBus_resp_data_3_data,
  output        io_dataWriteBus_req_valid,
  output [9:0]  io_dataWriteBus_req_bits_setIdx,
  output [63:0] io_dataWriteBus_req_bits_data_data,
  output [3:0]  io_dataWriteBus_req_bits_waymask,
  output        io_metaWriteBus_req_valid,
  output [6:0]  io_metaWriteBus_req_bits_setIdx,
  output [18:0] io_metaWriteBus_req_bits_data_tag,
  output        io_metaWriteBus_req_bits_data_valid,
  output        io_metaWriteBus_req_bits_data_dirty,
  output [3:0]  io_metaWriteBus_req_bits_waymask,
  input         io_mem_req_ready,
  output        io_mem_req_valid,
  output [31:0] io_mem_req_bits_addr,
  output [2:0]  io_mem_req_bits_size,
  output [3:0]  io_mem_req_bits_cmd,
  output [7:0]  io_mem_req_bits_wmask,
  output [63:0] io_mem_req_bits_wdata,
  output        io_mem_resp_ready,
  input         io_mem_resp_valid,
  input  [3:0]  io_mem_resp_bits_cmd,
  input  [63:0] io_mem_resp_bits_rdata,
  input         io_mmio_req_ready,
  output        io_mmio_req_valid,
  output [31:0] io_mmio_req_bits_addr,
  output        io_mmio_resp_ready,
  input         io_mmio_resp_valid,
  input  [63:0] io_mmio_resp_bits_rdata,
  output        io_cohResp_valid,
  input         DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
`endif // RANDOMIZE_REG_INIT
  wire  metaWriteArb_io_in_0_valid; // @[Cache.scala 241:28]
  wire [6:0] metaWriteArb_io_in_0_bits_setIdx; // @[Cache.scala 241:28]
  wire [18:0] metaWriteArb_io_in_0_bits_data_tag; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_in_0_bits_data_dirty; // @[Cache.scala 241:28]
  wire [3:0] metaWriteArb_io_in_0_bits_waymask; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_in_1_valid; // @[Cache.scala 241:28]
  wire [6:0] metaWriteArb_io_in_1_bits_setIdx; // @[Cache.scala 241:28]
  wire [18:0] metaWriteArb_io_in_1_bits_data_tag; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_in_1_bits_data_dirty; // @[Cache.scala 241:28]
  wire [3:0] metaWriteArb_io_in_1_bits_waymask; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_out_valid; // @[Cache.scala 241:28]
  wire [6:0] metaWriteArb_io_out_bits_setIdx; // @[Cache.scala 241:28]
  wire [18:0] metaWriteArb_io_out_bits_data_tag; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_out_bits_data_dirty; // @[Cache.scala 241:28]
  wire [3:0] metaWriteArb_io_out_bits_waymask; // @[Cache.scala 241:28]
  wire  dataWriteArb_io_in_0_valid; // @[Cache.scala 242:28]
  wire [9:0] dataWriteArb_io_in_0_bits_setIdx; // @[Cache.scala 242:28]
  wire [63:0] dataWriteArb_io_in_0_bits_data_data; // @[Cache.scala 242:28]
  wire [3:0] dataWriteArb_io_in_0_bits_waymask; // @[Cache.scala 242:28]
  wire  dataWriteArb_io_in_1_valid; // @[Cache.scala 242:28]
  wire [9:0] dataWriteArb_io_in_1_bits_setIdx; // @[Cache.scala 242:28]
  wire [63:0] dataWriteArb_io_in_1_bits_data_data; // @[Cache.scala 242:28]
  wire [3:0] dataWriteArb_io_in_1_bits_waymask; // @[Cache.scala 242:28]
  wire  dataWriteArb_io_out_valid; // @[Cache.scala 242:28]
  wire [9:0] dataWriteArb_io_out_bits_setIdx; // @[Cache.scala 242:28]
  wire [63:0] dataWriteArb_io_out_bits_data_data; // @[Cache.scala 242:28]
  wire [3:0] dataWriteArb_io_out_bits_waymask; // @[Cache.scala 242:28]
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[Cache.scala 245:31]
  wire [6:0] addr_index = io_in_bits_req_addr[12:6]; // @[Cache.scala 245:31]
  wire [18:0] addr_tag = io_in_bits_req_addr[31:13]; // @[Cache.scala 245:31]
  wire  mmio = io_in_valid & io_in_bits_mmio; // @[Cache.scala 246:26]
  wire  hit = io_in_valid & io_in_bits_hit; // @[Cache.scala 247:25]
  wire  _T_5 = ~io_in_bits_hit; // @[Cache.scala 248:29]
  wire  miss = io_in_valid & _T_5; // @[Cache.scala 248:26]
  wire [20:0] _T_14 = {io_in_bits_metas_0_tag,io_in_bits_metas_0_valid,io_in_bits_metas_0_dirty}; // @[Mux.scala 27:72]
  wire [20:0] _T_15 = io_in_bits_waymask[0] ? _T_14 : 21'h0; // @[Mux.scala 27:72]
  wire [20:0] _T_17 = {io_in_bits_metas_1_tag,io_in_bits_metas_1_valid,io_in_bits_metas_1_dirty}; // @[Mux.scala 27:72]
  wire [20:0] _T_18 = io_in_bits_waymask[1] ? _T_17 : 21'h0; // @[Mux.scala 27:72]
  wire [20:0] _T_20 = {io_in_bits_metas_2_tag,io_in_bits_metas_2_valid,io_in_bits_metas_2_dirty}; // @[Mux.scala 27:72]
  wire [20:0] _T_21 = io_in_bits_waymask[2] ? _T_20 : 21'h0; // @[Mux.scala 27:72]
  wire [20:0] _T_23 = {io_in_bits_metas_3_tag,io_in_bits_metas_3_valid,io_in_bits_metas_3_dirty}; // @[Mux.scala 27:72]
  wire [20:0] _T_24 = io_in_bits_waymask[3] ? _T_23 : 21'h0; // @[Mux.scala 27:72]
  wire [20:0] _T_25 = _T_15 | _T_18; // @[Mux.scala 27:72]
  wire [20:0] _T_26 = _T_25 | _T_21; // @[Mux.scala 27:72]
  wire [20:0] _T_27 = _T_26 | _T_24; // @[Mux.scala 27:72]
  wire [18:0] meta_tag = _T_27[20:2]; // @[Mux.scala 27:72]
  wire  _T_32 = mmio & hit; // @[Cache.scala 252:17]
  wire  _T_33 = ~_T_32; // @[Cache.scala 252:10]
  wire  _T_35 = _T_33 | reset; // @[Cache.scala 252:9]
  wire  _T_36 = ~_T_35; // @[Cache.scala 252:9]
  wire  _T_37 = io_in_bits_waymask == io_in_bits_forwardData_waymask; // @[Cache.scala 260:71]
  wire  useForwardData = io_in_bits_isForwardData & _T_37; // @[Cache.scala 260:49]
  wire [63:0] _T_42 = io_in_bits_waymask[0] ? io_in_bits_datas_0_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_43 = io_in_bits_waymask[1] ? io_in_bits_datas_1_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_44 = io_in_bits_waymask[2] ? io_in_bits_datas_2_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_45 = io_in_bits_waymask[3] ? io_in_bits_datas_3_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_46 = _T_42 | _T_43; // @[Mux.scala 27:72]
  wire [63:0] _T_47 = _T_46 | _T_44; // @[Mux.scala 27:72]
  wire [63:0] _T_48 = _T_47 | _T_45; // @[Mux.scala 27:72]
  wire [63:0] dataRead = useForwardData ? io_in_bits_forwardData_data_data : _T_48; // @[Cache.scala 262:21]
  wire  _T_86 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire [9:0] dataHitWriteBus_req_bits_setIdx = {addr_index,addr_wordIndex}; // @[Cat.scala 29:58]
  reg [3:0] state; // @[Cache.scala 281:22]
  reg  needFlush; // @[Cache.scala 282:26]
  wire  _T_114 = state != 4'h0; // @[Cache.scala 284:28]
  wire  _T_115 = io_flush & _T_114; // @[Cache.scala 284:18]
  wire  _GEN_1 = _T_115 | needFlush; // @[Cache.scala 284:41]
  wire  _T_117 = _T_86 & needFlush; // @[Cache.scala 285:23]
  reg [2:0] value_1; // @[Counter.scala 29:33]
  reg [2:0] value_2; // @[Counter.scala 29:33]
  reg [1:0] state2; // @[Cache.scala 291:23]
  wire  _T_118 = state == 4'h3; // @[Cache.scala 293:39]
  wire  _T_119 = state == 4'h8; // @[Cache.scala 293:66]
  wire  _T_120 = _T_118 | _T_119; // @[Cache.scala 293:57]
  wire  _T_121 = state2 == 2'h0; // @[Cache.scala 293:92]
  wire [2:0] _T_124 = _T_119 ? value_1 : value_2; // @[Cache.scala 294:33]
  wire  _T_126 = state2 == 2'h1; // @[Cache.scala 295:60]
  reg [63:0] dataWay_0_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_1_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_2_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_3_data; // @[Reg.scala 15:16]
  wire [63:0] _T_131 = io_in_bits_waymask[0] ? dataWay_0_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_132 = io_in_bits_waymask[1] ? dataWay_1_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_133 = io_in_bits_waymask[2] ? dataWay_2_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_134 = io_in_bits_waymask[3] ? dataWay_3_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_135 = _T_131 | _T_132; // @[Mux.scala 27:72]
  wire [63:0] _T_136 = _T_135 | _T_133; // @[Mux.scala 27:72]
  wire  _T_141 = 2'h0 == state2; // @[Conditional.scala 37:30]
  wire  _T_142 = io_dataReadBus_req_ready & io_dataReadBus_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_143 = 2'h1 == state2; // @[Conditional.scala 37:30]
  wire  _T_144 = 2'h2 == state2; // @[Conditional.scala 37:30]
  wire  _T_145 = io_mem_req_ready & io_mem_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_147 = _T_145 | io_cohResp_valid; // @[Cache.scala 301:46]
  wire [31:0] raddr = {io_in_bits_req_addr[31:3],3'h0}; // @[Cat.scala 29:58]
  wire [31:0] waddr = {meta_tag,addr_index,6'h0}; // @[Cat.scala 29:58]
  wire  _T_152 = state == 4'h1; // @[Cache.scala 309:23]
  wire  _T_153 = value_2 == 3'h7; // @[Cache.scala 310:29]
  wire [2:0] _T_154 = _T_153 ? 3'h7 : 3'h3; // @[Cache.scala 310:8]
  wire [2:0] cmd = _T_152 ? 3'h2 : _T_154; // @[Cache.scala 309:16]
  wire  _T_160 = state2 == 2'h2; // @[Cache.scala 316:89]
  wire  _T_161 = _T_118 & _T_160; // @[Cache.scala 316:78]
  reg  afterFirstRead; // @[Cache.scala 323:31]
  reg  alreadyOutFire; // @[Reg.scala 27:20]
  wire  _GEN_12 = _T_86 | alreadyOutFire; // @[Reg.scala 28:19]
  wire  _T_165 = ~afterFirstRead; // @[Cache.scala 325:22]
  wire  _T_166 = io_mem_resp_ready & io_mem_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_167 = _T_165 & _T_166; // @[Cache.scala 325:38]
  wire  _T_168 = state == 4'h2; // @[Cache.scala 325:70]
  wire  readingFirst = _T_167 & _T_168; // @[Cache.scala 325:60]
  wire  _T_170 = state == 4'h6; // @[Cache.scala 327:52]
  wire  _T_171 = mmio ? _T_170 : readingFirst; // @[Cache.scala 327:39]
  reg [63:0] inRdataRegDemand; // @[Reg.scala 15:16]
  wire  _T_172 = state == 4'h0; // @[Cache.scala 330:31]
  wire  _T_202 = 4'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_210 = miss | mmio; // @[Cache.scala 353:26]
  wire  _T_211 = ~io_flush; // @[Cache.scala 353:38]
  wire  _T_212 = _T_210 & _T_211; // @[Cache.scala 353:35]
  wire  _T_217 = 4'h5 == state; // @[Conditional.scala 37:30]
  wire  _T_218 = io_mmio_req_ready & io_mmio_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_219 = 4'h6 == state; // @[Conditional.scala 37:30]
  wire  _T_220 = io_mmio_resp_ready & io_mmio_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_221 = 4'h8 == state; // @[Conditional.scala 37:30]
  wire [2:0] _T_226 = value_1 + 3'h1; // @[Counter.scala 39:22]
  wire  _T_232 = 4'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_234 = 4'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_240 = io_mem_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire  _GEN_33 = _T_166 | afterFirstRead; // @[Cache.scala 372:33]
  wire  _T_241 = 4'h3 == state; // @[Conditional.scala 37:30]
  wire [2:0] _T_245 = value_2 + 3'h1; // @[Counter.scala 39:22]
  wire  _T_246 = io_mem_req_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_248 = _T_246 & _T_145; // @[Cache.scala 382:43]
  wire  _T_249 = 4'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_251 = 4'h7 == state; // @[Conditional.scala 37:30]
  wire  _T_253 = _T_86 | needFlush; // @[Cache.scala 386:44]
  wire  _T_254 = _T_253 | alreadyOutFire; // @[Cache.scala 386:57]
  wire  dataRefillWriteBus_req_valid = _T_168 & _T_166; // @[Cache.scala 391:39]
  wire  _T_293 = state == 4'h7; // @[Cache.scala 433:48]
  wire  _T_310 = ~alreadyOutFire; // @[Cache.scala 434:110]
  wire  _T_311 = afterFirstRead & _T_310; // @[Cache.scala 434:107]
  wire  _T_312 = mmio ? _T_293 : _T_311; // @[Cache.scala 434:45]
  wire  _T_313 = hit | _T_312; // @[Cache.scala 434:28]
  wire  _T_329 = _T_293 & _GEN_12; // @[Cache.scala 442:70]
  wire  _T_335 = io_out_ready & _T_172; // @[Cache.scala 445:31]
  wire  _T_336 = ~miss; // @[Cache.scala 445:73]
  wire [255:0] _T_371 = {io_in_bits_datas_3_data,io_in_bits_datas_2_data,io_in_bits_datas_1_data,io_in_bits_datas_0_data}; // @[Cache.scala 451:465]
  reg [63:0] _T_372; // @[GTimer.scala 24:20]
  wire [63:0] _T_374 = _T_372 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_378 = ~reset; // @[Debug.scala 56:24]
  reg [63:0] _T_382; // @[GTimer.scala 24:20]
  wire [63:0] _T_384 = _T_382 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_385; // @[GTimer.scala 24:20]
  wire [63:0] _T_387 = _T_385 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_389 = io_metaWriteBus_req_valid & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  reg [63:0] _T_394; // @[GTimer.scala 24:20]
  wire [63:0] _T_396 = _T_394 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_403; // @[GTimer.scala 24:20]
  wire [63:0] _T_405 = _T_403 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_412; // @[GTimer.scala 24:20]
  wire [63:0] _T_414 = _T_412 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_424; // @[GTimer.scala 24:20]
  wire [63:0] _T_426 = _T_424 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_433; // @[GTimer.scala 24:20]
  wire [63:0] _T_435 = _T_433 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_443; // @[GTimer.scala 24:20]
  wire [63:0] _T_445 = _T_443 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_447 = io_dataWriteBus_req_valid & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  wire  _T_454 = _T_118 & _T_145; // @[Cache.scala 460:35]
  reg [63:0] _T_461; // @[GTimer.scala 24:20]
  wire [63:0] _T_463 = _T_461 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_465 = _T_454 & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  wire  _T_472 = _T_152 & _T_145; // @[Cache.scala 461:34]
  reg [63:0] _T_479; // @[GTimer.scala 24:20]
  wire [63:0] _T_481 = _T_479 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_483 = _T_472 & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  reg [63:0] _T_497; // @[GTimer.scala 24:20]
  wire [63:0] _T_499 = _T_497 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_501 = dataRefillWriteBus_req_valid & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  Arbiter metaWriteArb ( // @[Cache.scala 241:28]
    .io_in_0_valid(metaWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(metaWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_tag(metaWriteArb_io_in_0_bits_data_tag),
    .io_in_0_bits_data_dirty(metaWriteArb_io_in_0_bits_data_dirty),
    .io_in_0_bits_waymask(metaWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(metaWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(metaWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_tag(metaWriteArb_io_in_1_bits_data_tag),
    .io_in_1_bits_data_dirty(metaWriteArb_io_in_1_bits_data_dirty),
    .io_in_1_bits_waymask(metaWriteArb_io_in_1_bits_waymask),
    .io_out_valid(metaWriteArb_io_out_valid),
    .io_out_bits_setIdx(metaWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_tag(metaWriteArb_io_out_bits_data_tag),
    .io_out_bits_data_dirty(metaWriteArb_io_out_bits_data_dirty),
    .io_out_bits_waymask(metaWriteArb_io_out_bits_waymask)
  );
  Arbiter_1 dataWriteArb ( // @[Cache.scala 242:28]
    .io_in_0_valid(dataWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(dataWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_data(dataWriteArb_io_in_0_bits_data_data),
    .io_in_0_bits_waymask(dataWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(dataWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(dataWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_data(dataWriteArb_io_in_1_bits_data_data),
    .io_in_1_bits_waymask(dataWriteArb_io_in_1_bits_waymask),
    .io_out_valid(dataWriteArb_io_out_valid),
    .io_out_bits_setIdx(dataWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_data(dataWriteArb_io_out_bits_data_data),
    .io_out_bits_waymask(dataWriteArb_io_out_bits_waymask)
  );
  assign io_in_ready = _T_335 & _T_336; // @[Cache.scala 445:15]
  assign io_out_valid = io_in_valid & _T_313; // @[Cache.scala 432:16]
  assign io_out_bits_cmd = 4'h6; // @[Cache.scala 427:21]
  assign io_out_bits_rdata = hit ? dataRead : inRdataRegDemand; // @[Cache.scala 426:23]
  assign io_out_bits_user = io_in_bits_req_user; // @[Cache.scala 429:56]
  assign io_isFinish = hit ? _T_86 : _T_329; // @[Cache.scala 441:15]
  assign io_dataReadBus_req_valid = _T_120 & _T_121; // @[SRAMTemplate.scala 53:20]
  assign io_dataReadBus_req_bits_setIdx = {addr_index,_T_124}; // @[SRAMTemplate.scala 26:17]
  assign io_dataWriteBus_req_valid = dataWriteArb_io_out_valid; // @[Cache.scala 396:23]
  assign io_dataWriteBus_req_bits_setIdx = dataWriteArb_io_out_bits_setIdx; // @[Cache.scala 396:23]
  assign io_dataWriteBus_req_bits_data_data = dataWriteArb_io_out_bits_data_data; // @[Cache.scala 396:23]
  assign io_dataWriteBus_req_bits_waymask = dataWriteArb_io_out_bits_waymask; // @[Cache.scala 396:23]
  assign io_metaWriteBus_req_valid = metaWriteArb_io_out_valid; // @[Cache.scala 406:23]
  assign io_metaWriteBus_req_bits_setIdx = metaWriteArb_io_out_bits_setIdx; // @[Cache.scala 406:23]
  assign io_metaWriteBus_req_bits_data_tag = metaWriteArb_io_out_bits_data_tag; // @[Cache.scala 406:23]
  assign io_metaWriteBus_req_bits_data_valid = 1'h1; // @[Cache.scala 406:23]
  assign io_metaWriteBus_req_bits_data_dirty = metaWriteArb_io_out_bits_data_dirty; // @[Cache.scala 406:23]
  assign io_metaWriteBus_req_bits_waymask = metaWriteArb_io_out_bits_waymask; // @[Cache.scala 406:23]
  assign io_mem_req_valid = _T_152 | _T_161; // @[Cache.scala 316:20]
  assign io_mem_req_bits_addr = _T_152 ? raddr : waddr; // @[SimpleBus.scala 64:15]
  assign io_mem_req_bits_size = 3'h3; // @[SimpleBus.scala 66:15]
  assign io_mem_req_bits_cmd = {{1'd0}, cmd}; // @[SimpleBus.scala 65:14]
  assign io_mem_req_bits_wmask = 8'hff; // @[SimpleBus.scala 68:16]
  assign io_mem_req_bits_wdata = _T_136 | _T_134; // @[SimpleBus.scala 67:16]
  assign io_mem_resp_ready = 1'h1; // @[Cache.scala 315:21]
  assign io_mmio_req_valid = state == 4'h5; // @[Cache.scala 321:21]
  assign io_mmio_req_bits_addr = io_in_bits_req_addr; // @[Cache.scala 319:20]
  assign io_mmio_resp_ready = 1'h1; // @[Cache.scala 320:22]
  assign io_cohResp_valid = _T_119 & _T_160; // @[Cache.scala 330:20]
  assign metaWriteArb_io_in_0_valid = 1'h0; // @[Cache.scala 404:25]
  assign metaWriteArb_io_in_0_bits_setIdx = io_in_bits_req_addr[12:6]; // @[Cache.scala 404:25]
  assign metaWriteArb_io_in_0_bits_data_tag = _T_27[20:2]; // @[Cache.scala 404:25]
  assign metaWriteArb_io_in_0_bits_data_dirty = 1'h0; // @[Cache.scala 404:25]
  assign metaWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[Cache.scala 404:25]
  assign metaWriteArb_io_in_1_valid = dataRefillWriteBus_req_valid & _T_240; // @[Cache.scala 405:25]
  assign metaWriteArb_io_in_1_bits_setIdx = io_in_bits_req_addr[12:6]; // @[Cache.scala 405:25]
  assign metaWriteArb_io_in_1_bits_data_tag = io_in_bits_req_addr[31:13]; // @[Cache.scala 405:25]
  assign metaWriteArb_io_in_1_bits_data_dirty = 1'h0; // @[Cache.scala 405:25]
  assign metaWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[Cache.scala 405:25]
  assign dataWriteArb_io_in_0_valid = 1'h0; // @[Cache.scala 394:25]
  assign dataWriteArb_io_in_0_bits_setIdx = {addr_index,addr_wordIndex}; // @[Cache.scala 394:25]
  assign dataWriteArb_io_in_0_bits_data_data = useForwardData ? io_in_bits_forwardData_data_data : _T_48; // @[Cache.scala 394:25]
  assign dataWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[Cache.scala 394:25]
  assign dataWriteArb_io_in_1_valid = _T_168 & _T_166; // @[Cache.scala 395:25]
  assign dataWriteArb_io_in_1_bits_setIdx = {addr_index,value_1}; // @[Cache.scala 395:25]
  assign dataWriteArb_io_in_1_bits_data_data = io_mem_resp_bits_rdata; // @[Cache.scala 395:25]
  assign dataWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[Cache.scala 395:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  needFlush = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  value_2 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  state2 = _RAND_4[1:0];
  _RAND_5 = {2{`RANDOM}};
  dataWay_0_data = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  dataWay_1_data = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  dataWay_2_data = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  dataWay_3_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  afterFirstRead = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  alreadyOutFire = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  inRdataRegDemand = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  _T_372 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  _T_382 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  _T_385 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  _T_394 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  _T_403 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  _T_412 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  _T_424 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  _T_433 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  _T_443 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  _T_461 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  _T_479 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  _T_497 = _RAND_23[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 4'h0;
    end else if (_T_202) begin
      if (_T_212) begin
        if (mmio) begin
          state <= 4'h5;
        end else begin
          state <= 4'h1;
        end
      end
    end else if (_T_217) begin
      if (_T_218) begin
        state <= 4'h6;
      end
    end else if (_T_219) begin
      if (_T_220) begin
        state <= 4'h7;
      end
    end else if (!(_T_221)) begin
      if (_T_232) begin
        if (_T_145) begin
          state <= 4'h2;
        end
      end else if (_T_234) begin
        if (_T_166) begin
          if (_T_240) begin
            state <= 4'h7;
          end
        end
      end else if (_T_241) begin
        if (_T_248) begin
          state <= 4'h4;
        end
      end else if (_T_249) begin
        if (_T_166) begin
          state <= 4'h1;
        end
      end else if (_T_251) begin
        if (_T_254) begin
          state <= 4'h0;
        end
      end
    end
    if (reset) begin
      needFlush <= 1'h0;
    end else if (_T_117) begin
      needFlush <= 1'h0;
    end else begin
      needFlush <= _GEN_1;
    end
    if (reset) begin
      value_1 <= 3'h0;
    end else if (!(_T_202)) begin
      if (!(_T_217)) begin
        if (!(_T_219)) begin
          if (_T_221) begin
            if (io_cohResp_valid) begin
              value_1 <= _T_226;
            end
          end else if (_T_232) begin
            if (_T_145) begin
              value_1 <= addr_wordIndex;
            end
          end else if (_T_234) begin
            if (_T_166) begin
              value_1 <= _T_226;
            end
          end
        end
      end
    end
    if (reset) begin
      value_2 <= 3'h0;
    end else if (!(_T_202)) begin
      if (!(_T_217)) begin
        if (!(_T_219)) begin
          if (!(_T_221)) begin
            if (!(_T_232)) begin
              if (!(_T_234)) begin
                if (_T_241) begin
                  if (_T_145) begin
                    value_2 <= _T_245;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      state2 <= 2'h0;
    end else if (_T_141) begin
      if (_T_142) begin
        state2 <= 2'h1;
      end
    end else if (_T_143) begin
      state2 <= 2'h2;
    end else if (_T_144) begin
      if (_T_147) begin
        state2 <= 2'h0;
      end
    end
    if (_T_126) begin
      dataWay_0_data <= io_dataReadBus_resp_data_0_data;
    end
    if (_T_126) begin
      dataWay_1_data <= io_dataReadBus_resp_data_1_data;
    end
    if (_T_126) begin
      dataWay_2_data <= io_dataReadBus_resp_data_2_data;
    end
    if (_T_126) begin
      dataWay_3_data <= io_dataReadBus_resp_data_3_data;
    end
    if (reset) begin
      afterFirstRead <= 1'h0;
    end else if (_T_202) begin
      afterFirstRead <= 1'h0;
    end else if (!(_T_217)) begin
      if (!(_T_219)) begin
        if (!(_T_221)) begin
          if (!(_T_232)) begin
            if (_T_234) begin
              afterFirstRead <= _GEN_33;
            end
          end
        end
      end
    end
    if (reset) begin
      alreadyOutFire <= 1'h0;
    end else if (_T_202) begin
      alreadyOutFire <= 1'h0;
    end else begin
      alreadyOutFire <= _GEN_12;
    end
    if (_T_171) begin
      if (mmio) begin
        inRdataRegDemand <= io_mmio_resp_bits_rdata;
      end else begin
        inRdataRegDemand <= io_mem_resp_bits_rdata;
      end
    end
    if (reset) begin
      _T_372 <= 64'h0;
    end else begin
      _T_372 <= _T_374;
    end
    if (reset) begin
      _T_382 <= 64'h0;
    end else begin
      _T_382 <= _T_384;
    end
    if (reset) begin
      _T_385 <= 64'h0;
    end else begin
      _T_385 <= _T_387;
    end
    if (reset) begin
      _T_394 <= 64'h0;
    end else begin
      _T_394 <= _T_396;
    end
    if (reset) begin
      _T_403 <= 64'h0;
    end else begin
      _T_403 <= _T_405;
    end
    if (reset) begin
      _T_412 <= 64'h0;
    end else begin
      _T_412 <= _T_414;
    end
    if (reset) begin
      _T_424 <= 64'h0;
    end else begin
      _T_424 <= _T_426;
    end
    if (reset) begin
      _T_433 <= 64'h0;
    end else begin
      _T_433 <= _T_435;
    end
    if (reset) begin
      _T_443 <= 64'h0;
    end else begin
      _T_443 <= _T_445;
    end
    if (reset) begin
      _T_461 <= 64'h0;
    end else begin
      _T_461 <= _T_463;
    end
    if (reset) begin
      _T_479 <= 64'h0;
    end else begin
      _T_479 <= _T_481;
    end
    if (reset) begin
      _T_497 <= 64'h0;
    end else begin
      _T_497 <= _T_499;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_36) begin
          $fwrite(32'h80000002,"Assertion failed: MMIO request should not hit in cache\n    at Cache.scala:252 assert(!(mmio && hit), \"MMIO request should not hit in cache\")\n"); // @[Cache.scala 252:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_36) begin
          $fatal; // @[Cache.scala 252:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_378) begin
          $fwrite(32'h80000002,"[%d] CacheStage3: ",_T_372); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_378) begin
          $fwrite(32'h80000002," metaread idx %x waymask %b metas %x%x:%x %x%x:%x %x%x:%x %x%x:%x %x\n",addr_index,io_in_bits_waymask,io_in_bits_metas_0_valid,io_in_bits_metas_0_dirty,io_in_bits_metas_0_tag,io_in_bits_metas_1_valid,io_in_bits_metas_1_dirty,io_in_bits_metas_1_tag,io_in_bits_metas_2_valid,io_in_bits_metas_2_dirty,io_in_bits_metas_2_tag,io_in_bits_metas_3_valid,io_in_bits_metas_3_dirty,io_in_bits_metas_3_tag,_T_371); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_389 & _T_378) begin
          $fwrite(32'h80000002,"[%d] CacheStage3: ",_T_385); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_389 & _T_378) begin
          $fwrite(32'h80000002,"%d: [icache S3]: metawrite idx %x wmask %b meta %x%x:%x\n",_T_382,io_metaWriteBus_req_bits_setIdx,io_metaWriteBus_req_bits_waymask,io_metaWriteBus_req_bits_data_valid,io_metaWriteBus_req_bits_data_dirty,io_metaWriteBus_req_bits_data_tag); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_378) begin
          $fwrite(32'h80000002,"[%d] CacheStage3: ",_T_394); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_378) begin
          $fwrite(32'h80000002," in.ready = %d, in.valid = %d, hit = %x, state = %d, addr = %x cmd:%d probe:%d isFinish:%d\n",io_in_ready,io_in_valid,hit,state,io_in_bits_req_addr,4'h0,1'h0,io_isFinish); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_378) begin
          $fwrite(32'h80000002,"[%d] CacheStage3: ",_T_403); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_378) begin
          $fwrite(32'h80000002," out.valid:%d rdata:%x cmd:%d user:%x id:%x \n",io_out_valid,io_out_bits_rdata,io_out_bits_cmd,io_out_bits_user,1'h0); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_378) begin
          $fwrite(32'h80000002,"[%d] CacheStage3: ",_T_412); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_378) begin
          $fwrite(32'h80000002," DHW: (%d, %d), data:%x setIdx:%x MHW:(%d, %d)\n",1'h0,1'h1,dataRead,dataHitWriteBus_req_bits_setIdx,1'h0,1'h1); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_378) begin
          $fwrite(32'h80000002,"[%d] CacheStage3: ",_T_424); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_378) begin
          $fwrite(32'h80000002," DreadCache: %x \n",_T_371); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_378) begin
          $fwrite(32'h80000002,"[%d] CacheStage3: ",_T_433); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_378) begin
          $fwrite(32'h80000002," useFD:%d isFD:%d FD:%x DreadArray:%x dataRead:%x inwaymask:%x FDwaymask:%x \n",useForwardData,io_in_bits_isForwardData,io_in_bits_forwardData_data_data,_T_48,dataRead,io_in_bits_waymask,io_in_bits_forwardData_waymask); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_447 & _T_378) begin
          $fwrite(32'h80000002,"[%d] CacheStage3: ",_T_443); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_447 & _T_378) begin
          $fwrite(32'h80000002,"[WB] waymask: %b data:%x setIdx:%x\n",io_dataWriteBus_req_bits_waymask,io_dataWriteBus_req_bits_data_data,io_dataWriteBus_req_bits_setIdx); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_465 & _T_378) begin
          $fwrite(32'h80000002,"[%d] CacheStage3: ",_T_461); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_465 & _T_378) begin
          $fwrite(32'h80000002,"[COUTW] cnt %x addr %x data %x cmd %x size %x wmask %x tag %x idx %x waymask %b \n",value_2,io_mem_req_bits_addr,io_mem_req_bits_wdata,io_mem_req_bits_cmd,io_mem_req_bits_size,io_mem_req_bits_wmask,addr_tag,addr_index,io_in_bits_waymask); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_483 & _T_378) begin
          $fwrite(32'h80000002,"[%d] CacheStage3: ",_T_479); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_483 & _T_378) begin
          $fwrite(32'h80000002,"[COUTR] addr %x tag %x idx %x waymask %b \n",io_mem_req_bits_addr,addr_tag,addr_index,io_in_bits_waymask); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_501 & _T_378) begin
          $fwrite(32'h80000002,"[%d] CacheStage3: ",_T_497); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_501 & _T_378) begin
          $fwrite(32'h80000002,"[COUTR] cnt %x data %x tag %x idx %x waymask %b \n",value_1,io_mem_resp_bits_rdata,addr_tag,addr_index,io_in_bits_waymask); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module SRAMTemplate_1(
  input         clock,
  input         reset,
  output        io_r_req_ready,
  input         io_r_req_valid,
  input  [6:0]  io_r_req_bits_setIdx,
  output [18:0] io_r_resp_data_0_tag,
  output        io_r_resp_data_0_valid,
  output        io_r_resp_data_0_dirty,
  output [18:0] io_r_resp_data_1_tag,
  output        io_r_resp_data_1_valid,
  output        io_r_resp_data_1_dirty,
  output [18:0] io_r_resp_data_2_tag,
  output        io_r_resp_data_2_valid,
  output        io_r_resp_data_2_dirty,
  output [18:0] io_r_resp_data_3_tag,
  output        io_r_resp_data_3_valid,
  output        io_r_resp_data_3_dirty,
  input         io_w_req_valid,
  input  [6:0]  io_w_req_bits_setIdx,
  input  [18:0] io_w_req_bits_data_tag,
  input         io_w_req_bits_data_dirty,
  input  [3:0]  io_w_req_bits_waymask
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  reg [20:0] array_0 [0:127]; // @[SRAMTemplate.scala 76:26]
  wire [20:0] array_0__T_21_data; // @[SRAMTemplate.scala 76:26]
  wire [6:0] array_0__T_21_addr; // @[SRAMTemplate.scala 76:26]
  wire [20:0] array_0__T_17_data; // @[SRAMTemplate.scala 76:26]
  wire [6:0] array_0__T_17_addr; // @[SRAMTemplate.scala 76:26]
  wire  array_0__T_17_mask; // @[SRAMTemplate.scala 76:26]
  wire  array_0__T_17_en; // @[SRAMTemplate.scala 76:26]
  reg  array_0__T_21_en_pipe_0;
  reg [6:0] array_0__T_21_addr_pipe_0;
  reg [20:0] array_1 [0:127]; // @[SRAMTemplate.scala 76:26]
  wire [20:0] array_1__T_21_data; // @[SRAMTemplate.scala 76:26]
  wire [6:0] array_1__T_21_addr; // @[SRAMTemplate.scala 76:26]
  wire [20:0] array_1__T_17_data; // @[SRAMTemplate.scala 76:26]
  wire [6:0] array_1__T_17_addr; // @[SRAMTemplate.scala 76:26]
  wire  array_1__T_17_mask; // @[SRAMTemplate.scala 76:26]
  wire  array_1__T_17_en; // @[SRAMTemplate.scala 76:26]
  reg  array_1__T_21_en_pipe_0;
  reg [6:0] array_1__T_21_addr_pipe_0;
  reg [20:0] array_2 [0:127]; // @[SRAMTemplate.scala 76:26]
  wire [20:0] array_2__T_21_data; // @[SRAMTemplate.scala 76:26]
  wire [6:0] array_2__T_21_addr; // @[SRAMTemplate.scala 76:26]
  wire [20:0] array_2__T_17_data; // @[SRAMTemplate.scala 76:26]
  wire [6:0] array_2__T_17_addr; // @[SRAMTemplate.scala 76:26]
  wire  array_2__T_17_mask; // @[SRAMTemplate.scala 76:26]
  wire  array_2__T_17_en; // @[SRAMTemplate.scala 76:26]
  reg  array_2__T_21_en_pipe_0;
  reg [6:0] array_2__T_21_addr_pipe_0;
  reg [20:0] array_3 [0:127]; // @[SRAMTemplate.scala 76:26]
  wire [20:0] array_3__T_21_data; // @[SRAMTemplate.scala 76:26]
  wire [6:0] array_3__T_21_addr; // @[SRAMTemplate.scala 76:26]
  wire [20:0] array_3__T_17_data; // @[SRAMTemplate.scala 76:26]
  wire [6:0] array_3__T_17_addr; // @[SRAMTemplate.scala 76:26]
  wire  array_3__T_17_mask; // @[SRAMTemplate.scala 76:26]
  wire  array_3__T_17_en; // @[SRAMTemplate.scala 76:26]
  reg  array_3__T_21_en_pipe_0;
  reg [6:0] array_3__T_21_addr_pipe_0;
  reg  resetState; // @[SRAMTemplate.scala 80:30]
  reg [6:0] resetSet; // @[Counter.scala 29:33]
  wire  _T_3 = resetSet == 7'h7f; // @[Counter.scala 38:24]
  wire [6:0] _T_5 = resetSet + 7'h1; // @[Counter.scala 39:22]
  wire  _GEN_1 = resetState & _T_3; // @[Counter.scala 67:17]
  wire  _GEN_2 = _GEN_1 ? 1'h0 : resetState; // @[SRAMTemplate.scala 82:24]
  wire  wen = io_w_req_valid | resetState; // @[SRAMTemplate.scala 88:52]
  wire  _T_6 = ~wen; // @[SRAMTemplate.scala 89:41]
  wire [20:0] _T_9 = {io_w_req_bits_data_tag,1'h1,io_w_req_bits_data_dirty}; // @[SRAMTemplate.scala 92:78]
  wire [3:0] waymask = resetState ? 4'hf : io_w_req_bits_waymask; // @[SRAMTemplate.scala 93:20]
  wire [20:0] _T_22 = array_0__T_21_data;
  wire [20:0] _T_26 = array_1__T_21_data;
  wire [20:0] _T_30 = array_2__T_21_data;
  wire [20:0] _T_34 = array_3__T_21_data;
  wire  _T_39 = ~resetState; // @[SRAMTemplate.scala 101:21]
  assign array_0__T_21_addr = array_0__T_21_addr_pipe_0;
  assign array_0__T_21_data = array_0[array_0__T_21_addr]; // @[SRAMTemplate.scala 76:26]
  assign array_0__T_17_data = resetState ? 21'h0 : _T_9;
  assign array_0__T_17_addr = resetState ? resetSet : io_w_req_bits_setIdx;
  assign array_0__T_17_mask = waymask[0];
  assign array_0__T_17_en = io_w_req_valid | resetState;
  assign array_1__T_21_addr = array_1__T_21_addr_pipe_0;
  assign array_1__T_21_data = array_1[array_1__T_21_addr]; // @[SRAMTemplate.scala 76:26]
  assign array_1__T_17_data = resetState ? 21'h0 : _T_9;
  assign array_1__T_17_addr = resetState ? resetSet : io_w_req_bits_setIdx;
  assign array_1__T_17_mask = waymask[1];
  assign array_1__T_17_en = io_w_req_valid | resetState;
  assign array_2__T_21_addr = array_2__T_21_addr_pipe_0;
  assign array_2__T_21_data = array_2[array_2__T_21_addr]; // @[SRAMTemplate.scala 76:26]
  assign array_2__T_17_data = resetState ? 21'h0 : _T_9;
  assign array_2__T_17_addr = resetState ? resetSet : io_w_req_bits_setIdx;
  assign array_2__T_17_mask = waymask[2];
  assign array_2__T_17_en = io_w_req_valid | resetState;
  assign array_3__T_21_addr = array_3__T_21_addr_pipe_0;
  assign array_3__T_21_data = array_3[array_3__T_21_addr]; // @[SRAMTemplate.scala 76:26]
  assign array_3__T_17_data = resetState ? 21'h0 : _T_9;
  assign array_3__T_17_addr = resetState ? resetSet : io_w_req_bits_setIdx;
  assign array_3__T_17_mask = waymask[3];
  assign array_3__T_17_en = io_w_req_valid | resetState;
  assign io_r_req_ready = _T_39 & _T_6; // @[SRAMTemplate.scala 101:18]
  assign io_r_resp_data_0_tag = _T_22[20:2]; // @[SRAMTemplate.scala 99:18]
  assign io_r_resp_data_0_valid = _T_22[1]; // @[SRAMTemplate.scala 99:18]
  assign io_r_resp_data_0_dirty = _T_22[0]; // @[SRAMTemplate.scala 99:18]
  assign io_r_resp_data_1_tag = _T_26[20:2]; // @[SRAMTemplate.scala 99:18]
  assign io_r_resp_data_1_valid = _T_26[1]; // @[SRAMTemplate.scala 99:18]
  assign io_r_resp_data_1_dirty = _T_26[0]; // @[SRAMTemplate.scala 99:18]
  assign io_r_resp_data_2_tag = _T_30[20:2]; // @[SRAMTemplate.scala 99:18]
  assign io_r_resp_data_2_valid = _T_30[1]; // @[SRAMTemplate.scala 99:18]
  assign io_r_resp_data_2_dirty = _T_30[0]; // @[SRAMTemplate.scala 99:18]
  assign io_r_resp_data_3_tag = _T_34[20:2]; // @[SRAMTemplate.scala 99:18]
  assign io_r_resp_data_3_valid = _T_34[1]; // @[SRAMTemplate.scala 99:18]
  assign io_r_resp_data_3_dirty = _T_34[0]; // @[SRAMTemplate.scala 99:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    array_0[initvar] = _RAND_0[20:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    array_1[initvar] = _RAND_3[20:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    array_2[initvar] = _RAND_6[20:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    array_3[initvar] = _RAND_9[20:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  array_0__T_21_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  array_0__T_21_addr_pipe_0 = _RAND_2[6:0];
  _RAND_4 = {1{`RANDOM}};
  array_1__T_21_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  array_1__T_21_addr_pipe_0 = _RAND_5[6:0];
  _RAND_7 = {1{`RANDOM}};
  array_2__T_21_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  array_2__T_21_addr_pipe_0 = _RAND_8[6:0];
  _RAND_10 = {1{`RANDOM}};
  array_3__T_21_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  array_3__T_21_addr_pipe_0 = _RAND_11[6:0];
  _RAND_12 = {1{`RANDOM}};
  resetState = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  resetSet = _RAND_13[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(array_0__T_17_en & array_0__T_17_mask) begin
      array_0[array_0__T_17_addr] <= array_0__T_17_data; // @[SRAMTemplate.scala 76:26]
    end
    array_0__T_21_en_pipe_0 <= io_r_req_valid & _T_6;
    if (io_r_req_valid & _T_6) begin
      array_0__T_21_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if(array_1__T_17_en & array_1__T_17_mask) begin
      array_1[array_1__T_17_addr] <= array_1__T_17_data; // @[SRAMTemplate.scala 76:26]
    end
    array_1__T_21_en_pipe_0 <= io_r_req_valid & _T_6;
    if (io_r_req_valid & _T_6) begin
      array_1__T_21_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if(array_2__T_17_en & array_2__T_17_mask) begin
      array_2[array_2__T_17_addr] <= array_2__T_17_data; // @[SRAMTemplate.scala 76:26]
    end
    array_2__T_21_en_pipe_0 <= io_r_req_valid & _T_6;
    if (io_r_req_valid & _T_6) begin
      array_2__T_21_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if(array_3__T_17_en & array_3__T_17_mask) begin
      array_3[array_3__T_17_addr] <= array_3__T_17_data; // @[SRAMTemplate.scala 76:26]
    end
    array_3__T_21_en_pipe_0 <= io_r_req_valid & _T_6;
    if (io_r_req_valid & _T_6) begin
      array_3__T_21_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    resetState <= reset | _GEN_2;
    if (reset) begin
      resetSet <= 7'h0;
    end else if (resetState) begin
      resetSet <= _T_5;
    end
  end
endmodule
module Arbiter_2(
  output       io_in_0_ready,
  input        io_in_0_valid,
  input  [6:0] io_in_0_bits_setIdx,
  input        io_out_ready,
  output       io_out_valid,
  output [6:0] io_out_bits_setIdx
);
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:14]
  assign io_out_valid = io_in_0_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_setIdx = io_in_0_bits_setIdx; // @[Arbiter.scala 124:15]
endmodule
module SRAMTemplateWithArbiter(
  input         clock,
  input         reset,
  output        io_r_0_req_ready,
  input         io_r_0_req_valid,
  input  [6:0]  io_r_0_req_bits_setIdx,
  output [18:0] io_r_0_resp_data_0_tag,
  output        io_r_0_resp_data_0_valid,
  output        io_r_0_resp_data_0_dirty,
  output [18:0] io_r_0_resp_data_1_tag,
  output        io_r_0_resp_data_1_valid,
  output        io_r_0_resp_data_1_dirty,
  output [18:0] io_r_0_resp_data_2_tag,
  output        io_r_0_resp_data_2_valid,
  output        io_r_0_resp_data_2_dirty,
  output [18:0] io_r_0_resp_data_3_tag,
  output        io_r_0_resp_data_3_valid,
  output        io_r_0_resp_data_3_dirty,
  input         io_w_req_valid,
  input  [6:0]  io_w_req_bits_setIdx,
  input  [18:0] io_w_req_bits_data_tag,
  input         io_w_req_bits_data_dirty,
  input  [3:0]  io_w_req_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  ram_clock; // @[SRAMTemplate.scala 121:19]
  wire  ram_reset; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_r_req_ready; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_r_req_valid; // @[SRAMTemplate.scala 121:19]
  wire [6:0] ram_io_r_req_bits_setIdx; // @[SRAMTemplate.scala 121:19]
  wire [18:0] ram_io_r_resp_data_0_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_r_resp_data_0_valid; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_r_resp_data_0_dirty; // @[SRAMTemplate.scala 121:19]
  wire [18:0] ram_io_r_resp_data_1_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_r_resp_data_1_valid; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_r_resp_data_1_dirty; // @[SRAMTemplate.scala 121:19]
  wire [18:0] ram_io_r_resp_data_2_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_r_resp_data_2_valid; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_r_resp_data_2_dirty; // @[SRAMTemplate.scala 121:19]
  wire [18:0] ram_io_r_resp_data_3_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_r_resp_data_3_valid; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_r_resp_data_3_dirty; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_w_req_valid; // @[SRAMTemplate.scala 121:19]
  wire [6:0] ram_io_w_req_bits_setIdx; // @[SRAMTemplate.scala 121:19]
  wire [18:0] ram_io_w_req_bits_data_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_w_req_bits_data_dirty; // @[SRAMTemplate.scala 121:19]
  wire [3:0] ram_io_w_req_bits_waymask; // @[SRAMTemplate.scala 121:19]
  wire  readArb_io_in_0_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_in_0_valid; // @[SRAMTemplate.scala 124:23]
  wire [6:0] readArb_io_in_0_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_out_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_out_valid; // @[SRAMTemplate.scala 124:23]
  wire [6:0] readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  reg  _T_1; // @[SRAMTemplate.scala 130:58]
  reg [18:0] _T_3_0_tag; // @[Reg.scala 27:20]
  reg  _T_3_0_valid; // @[Reg.scala 27:20]
  reg  _T_3_0_dirty; // @[Reg.scala 27:20]
  reg [18:0] _T_3_1_tag; // @[Reg.scala 27:20]
  reg  _T_3_1_valid; // @[Reg.scala 27:20]
  reg  _T_3_1_dirty; // @[Reg.scala 27:20]
  reg [18:0] _T_3_2_tag; // @[Reg.scala 27:20]
  reg  _T_3_2_valid; // @[Reg.scala 27:20]
  reg  _T_3_2_dirty; // @[Reg.scala 27:20]
  reg [18:0] _T_3_3_tag; // @[Reg.scala 27:20]
  reg  _T_3_3_valid; // @[Reg.scala 27:20]
  reg  _T_3_3_dirty; // @[Reg.scala 27:20]
  SRAMTemplate_1 ram ( // @[SRAMTemplate.scala 121:19]
    .clock(ram_clock),
    .reset(ram_reset),
    .io_r_req_ready(ram_io_r_req_ready),
    .io_r_req_valid(ram_io_r_req_valid),
    .io_r_req_bits_setIdx(ram_io_r_req_bits_setIdx),
    .io_r_resp_data_0_tag(ram_io_r_resp_data_0_tag),
    .io_r_resp_data_0_valid(ram_io_r_resp_data_0_valid),
    .io_r_resp_data_0_dirty(ram_io_r_resp_data_0_dirty),
    .io_r_resp_data_1_tag(ram_io_r_resp_data_1_tag),
    .io_r_resp_data_1_valid(ram_io_r_resp_data_1_valid),
    .io_r_resp_data_1_dirty(ram_io_r_resp_data_1_dirty),
    .io_r_resp_data_2_tag(ram_io_r_resp_data_2_tag),
    .io_r_resp_data_2_valid(ram_io_r_resp_data_2_valid),
    .io_r_resp_data_2_dirty(ram_io_r_resp_data_2_dirty),
    .io_r_resp_data_3_tag(ram_io_r_resp_data_3_tag),
    .io_r_resp_data_3_valid(ram_io_r_resp_data_3_valid),
    .io_r_resp_data_3_dirty(ram_io_r_resp_data_3_dirty),
    .io_w_req_valid(ram_io_w_req_valid),
    .io_w_req_bits_setIdx(ram_io_w_req_bits_setIdx),
    .io_w_req_bits_data_tag(ram_io_w_req_bits_data_tag),
    .io_w_req_bits_data_dirty(ram_io_w_req_bits_data_dirty),
    .io_w_req_bits_waymask(ram_io_w_req_bits_waymask)
  );
  Arbiter_2 readArb ( // @[SRAMTemplate.scala 124:23]
    .io_in_0_ready(readArb_io_in_0_ready),
    .io_in_0_valid(readArb_io_in_0_valid),
    .io_in_0_bits_setIdx(readArb_io_in_0_bits_setIdx),
    .io_out_ready(readArb_io_out_ready),
    .io_out_valid(readArb_io_out_valid),
    .io_out_bits_setIdx(readArb_io_out_bits_setIdx)
  );
  assign io_r_0_req_ready = readArb_io_in_0_ready; // @[SRAMTemplate.scala 125:17]
  assign io_r_0_resp_data_0_tag = _T_1 ? ram_io_r_resp_data_0_tag : _T_3_0_tag; // @[SRAMTemplate.scala 130:17]
  assign io_r_0_resp_data_0_valid = _T_1 ? ram_io_r_resp_data_0_valid : _T_3_0_valid; // @[SRAMTemplate.scala 130:17]
  assign io_r_0_resp_data_0_dirty = _T_1 ? ram_io_r_resp_data_0_dirty : _T_3_0_dirty; // @[SRAMTemplate.scala 130:17]
  assign io_r_0_resp_data_1_tag = _T_1 ? ram_io_r_resp_data_1_tag : _T_3_1_tag; // @[SRAMTemplate.scala 130:17]
  assign io_r_0_resp_data_1_valid = _T_1 ? ram_io_r_resp_data_1_valid : _T_3_1_valid; // @[SRAMTemplate.scala 130:17]
  assign io_r_0_resp_data_1_dirty = _T_1 ? ram_io_r_resp_data_1_dirty : _T_3_1_dirty; // @[SRAMTemplate.scala 130:17]
  assign io_r_0_resp_data_2_tag = _T_1 ? ram_io_r_resp_data_2_tag : _T_3_2_tag; // @[SRAMTemplate.scala 130:17]
  assign io_r_0_resp_data_2_valid = _T_1 ? ram_io_r_resp_data_2_valid : _T_3_2_valid; // @[SRAMTemplate.scala 130:17]
  assign io_r_0_resp_data_2_dirty = _T_1 ? ram_io_r_resp_data_2_dirty : _T_3_2_dirty; // @[SRAMTemplate.scala 130:17]
  assign io_r_0_resp_data_3_tag = _T_1 ? ram_io_r_resp_data_3_tag : _T_3_3_tag; // @[SRAMTemplate.scala 130:17]
  assign io_r_0_resp_data_3_valid = _T_1 ? ram_io_r_resp_data_3_valid : _T_3_3_valid; // @[SRAMTemplate.scala 130:17]
  assign io_r_0_resp_data_3_dirty = _T_1 ? ram_io_r_resp_data_3_dirty : _T_3_3_dirty; // @[SRAMTemplate.scala 130:17]
  assign ram_clock = clock;
  assign ram_reset = reset;
  assign ram_io_r_req_valid = readArb_io_out_valid; // @[SRAMTemplate.scala 126:16]
  assign ram_io_r_req_bits_setIdx = readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 126:16]
  assign ram_io_w_req_valid = io_w_req_valid; // @[SRAMTemplate.scala 122:12]
  assign ram_io_w_req_bits_setIdx = io_w_req_bits_setIdx; // @[SRAMTemplate.scala 122:12]
  assign ram_io_w_req_bits_data_tag = io_w_req_bits_data_tag; // @[SRAMTemplate.scala 122:12]
  assign ram_io_w_req_bits_data_dirty = io_w_req_bits_data_dirty; // @[SRAMTemplate.scala 122:12]
  assign ram_io_w_req_bits_waymask = io_w_req_bits_waymask; // @[SRAMTemplate.scala 122:12]
  assign readArb_io_in_0_valid = io_r_0_req_valid; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_in_0_bits_setIdx = io_r_0_req_bits_setIdx; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_out_ready = ram_io_r_req_ready; // @[SRAMTemplate.scala 126:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _T_3_0_tag = _RAND_1[18:0];
  _RAND_2 = {1{`RANDOM}};
  _T_3_0_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _T_3_0_dirty = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_3_1_tag = _RAND_4[18:0];
  _RAND_5 = {1{`RANDOM}};
  _T_3_1_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _T_3_1_dirty = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_3_2_tag = _RAND_7[18:0];
  _RAND_8 = {1{`RANDOM}};
  _T_3_2_valid = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _T_3_2_dirty = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _T_3_3_tag = _RAND_10[18:0];
  _RAND_11 = {1{`RANDOM}};
  _T_3_3_valid = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _T_3_3_dirty = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_1 <= io_r_0_req_ready & io_r_0_req_valid;
    if (reset) begin
      _T_3_0_tag <= 19'h0;
    end else if (_T_1) begin
      _T_3_0_tag <= ram_io_r_resp_data_0_tag;
    end
    if (reset) begin
      _T_3_0_valid <= 1'h0;
    end else if (_T_1) begin
      _T_3_0_valid <= ram_io_r_resp_data_0_valid;
    end
    if (reset) begin
      _T_3_0_dirty <= 1'h0;
    end else if (_T_1) begin
      _T_3_0_dirty <= ram_io_r_resp_data_0_dirty;
    end
    if (reset) begin
      _T_3_1_tag <= 19'h0;
    end else if (_T_1) begin
      _T_3_1_tag <= ram_io_r_resp_data_1_tag;
    end
    if (reset) begin
      _T_3_1_valid <= 1'h0;
    end else if (_T_1) begin
      _T_3_1_valid <= ram_io_r_resp_data_1_valid;
    end
    if (reset) begin
      _T_3_1_dirty <= 1'h0;
    end else if (_T_1) begin
      _T_3_1_dirty <= ram_io_r_resp_data_1_dirty;
    end
    if (reset) begin
      _T_3_2_tag <= 19'h0;
    end else if (_T_1) begin
      _T_3_2_tag <= ram_io_r_resp_data_2_tag;
    end
    if (reset) begin
      _T_3_2_valid <= 1'h0;
    end else if (_T_1) begin
      _T_3_2_valid <= ram_io_r_resp_data_2_valid;
    end
    if (reset) begin
      _T_3_2_dirty <= 1'h0;
    end else if (_T_1) begin
      _T_3_2_dirty <= ram_io_r_resp_data_2_dirty;
    end
    if (reset) begin
      _T_3_3_tag <= 19'h0;
    end else if (_T_1) begin
      _T_3_3_tag <= ram_io_r_resp_data_3_tag;
    end
    if (reset) begin
      _T_3_3_valid <= 1'h0;
    end else if (_T_1) begin
      _T_3_3_valid <= ram_io_r_resp_data_3_valid;
    end
    if (reset) begin
      _T_3_3_dirty <= 1'h0;
    end else if (_T_1) begin
      _T_3_3_dirty <= ram_io_r_resp_data_3_dirty;
    end
  end
endmodule
module SRAMTemplate_2(
  input         clock,
  output        io_r_req_ready,
  input         io_r_req_valid,
  input  [9:0]  io_r_req_bits_setIdx,
  output [63:0] io_r_resp_data_0_data,
  output [63:0] io_r_resp_data_1_data,
  output [63:0] io_r_resp_data_2_data,
  output [63:0] io_r_resp_data_3_data,
  input         io_w_req_valid,
  input  [9:0]  io_w_req_bits_setIdx,
  input  [63:0] io_w_req_bits_data_data,
  input  [3:0]  io_w_req_bits_waymask
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_9;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] array_0 [0:1023]; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_0__T_13_data; // @[SRAMTemplate.scala 76:26]
  wire [9:0] array_0__T_13_addr; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_0__T_9_data; // @[SRAMTemplate.scala 76:26]
  wire [9:0] array_0__T_9_addr; // @[SRAMTemplate.scala 76:26]
  wire  array_0__T_9_mask; // @[SRAMTemplate.scala 76:26]
  wire  array_0__T_9_en; // @[SRAMTemplate.scala 76:26]
  reg  array_0__T_13_en_pipe_0;
  reg [9:0] array_0__T_13_addr_pipe_0;
  reg [63:0] array_1 [0:1023]; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_1__T_13_data; // @[SRAMTemplate.scala 76:26]
  wire [9:0] array_1__T_13_addr; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_1__T_9_data; // @[SRAMTemplate.scala 76:26]
  wire [9:0] array_1__T_9_addr; // @[SRAMTemplate.scala 76:26]
  wire  array_1__T_9_mask; // @[SRAMTemplate.scala 76:26]
  wire  array_1__T_9_en; // @[SRAMTemplate.scala 76:26]
  reg  array_1__T_13_en_pipe_0;
  reg [9:0] array_1__T_13_addr_pipe_0;
  reg [63:0] array_2 [0:1023]; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_2__T_13_data; // @[SRAMTemplate.scala 76:26]
  wire [9:0] array_2__T_13_addr; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_2__T_9_data; // @[SRAMTemplate.scala 76:26]
  wire [9:0] array_2__T_9_addr; // @[SRAMTemplate.scala 76:26]
  wire  array_2__T_9_mask; // @[SRAMTemplate.scala 76:26]
  wire  array_2__T_9_en; // @[SRAMTemplate.scala 76:26]
  reg  array_2__T_13_en_pipe_0;
  reg [9:0] array_2__T_13_addr_pipe_0;
  reg [63:0] array_3 [0:1023]; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_3__T_13_data; // @[SRAMTemplate.scala 76:26]
  wire [9:0] array_3__T_13_addr; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_3__T_9_data; // @[SRAMTemplate.scala 76:26]
  wire [9:0] array_3__T_9_addr; // @[SRAMTemplate.scala 76:26]
  wire  array_3__T_9_mask; // @[SRAMTemplate.scala 76:26]
  wire  array_3__T_9_en; // @[SRAMTemplate.scala 76:26]
  reg  array_3__T_13_en_pipe_0;
  reg [9:0] array_3__T_13_addr_pipe_0;
  wire  _T = ~io_w_req_valid; // @[SRAMTemplate.scala 89:41]
  assign array_0__T_13_addr = array_0__T_13_addr_pipe_0;
  assign array_0__T_13_data = array_0[array_0__T_13_addr]; // @[SRAMTemplate.scala 76:26]
  assign array_0__T_9_data = io_w_req_bits_data_data;
  assign array_0__T_9_addr = io_w_req_bits_setIdx;
  assign array_0__T_9_mask = io_w_req_bits_waymask[0];
  assign array_0__T_9_en = io_w_req_valid;
  assign array_1__T_13_addr = array_1__T_13_addr_pipe_0;
  assign array_1__T_13_data = array_1[array_1__T_13_addr]; // @[SRAMTemplate.scala 76:26]
  assign array_1__T_9_data = io_w_req_bits_data_data;
  assign array_1__T_9_addr = io_w_req_bits_setIdx;
  assign array_1__T_9_mask = io_w_req_bits_waymask[1];
  assign array_1__T_9_en = io_w_req_valid;
  assign array_2__T_13_addr = array_2__T_13_addr_pipe_0;
  assign array_2__T_13_data = array_2[array_2__T_13_addr]; // @[SRAMTemplate.scala 76:26]
  assign array_2__T_9_data = io_w_req_bits_data_data;
  assign array_2__T_9_addr = io_w_req_bits_setIdx;
  assign array_2__T_9_mask = io_w_req_bits_waymask[2];
  assign array_2__T_9_en = io_w_req_valid;
  assign array_3__T_13_addr = array_3__T_13_addr_pipe_0;
  assign array_3__T_13_data = array_3[array_3__T_13_addr]; // @[SRAMTemplate.scala 76:26]
  assign array_3__T_9_data = io_w_req_bits_data_data;
  assign array_3__T_9_addr = io_w_req_bits_setIdx;
  assign array_3__T_9_mask = io_w_req_bits_waymask[3];
  assign array_3__T_9_en = io_w_req_valid;
  assign io_r_req_ready = ~io_w_req_valid; // @[SRAMTemplate.scala 101:18]
  assign io_r_resp_data_0_data = array_0__T_13_data; // @[SRAMTemplate.scala 99:18]
  assign io_r_resp_data_1_data = array_1__T_13_data; // @[SRAMTemplate.scala 99:18]
  assign io_r_resp_data_2_data = array_2__T_13_data; // @[SRAMTemplate.scala 99:18]
  assign io_r_resp_data_3_data = array_3__T_13_data; // @[SRAMTemplate.scala 99:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    array_0[initvar] = _RAND_0[63:0];
  _RAND_3 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    array_1[initvar] = _RAND_3[63:0];
  _RAND_6 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    array_2[initvar] = _RAND_6[63:0];
  _RAND_9 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    array_3[initvar] = _RAND_9[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  array_0__T_13_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  array_0__T_13_addr_pipe_0 = _RAND_2[9:0];
  _RAND_4 = {1{`RANDOM}};
  array_1__T_13_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  array_1__T_13_addr_pipe_0 = _RAND_5[9:0];
  _RAND_7 = {1{`RANDOM}};
  array_2__T_13_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  array_2__T_13_addr_pipe_0 = _RAND_8[9:0];
  _RAND_10 = {1{`RANDOM}};
  array_3__T_13_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  array_3__T_13_addr_pipe_0 = _RAND_11[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(array_0__T_9_en & array_0__T_9_mask) begin
      array_0[array_0__T_9_addr] <= array_0__T_9_data; // @[SRAMTemplate.scala 76:26]
    end
    array_0__T_13_en_pipe_0 <= io_r_req_valid & _T;
    if (io_r_req_valid & _T) begin
      array_0__T_13_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if(array_1__T_9_en & array_1__T_9_mask) begin
      array_1[array_1__T_9_addr] <= array_1__T_9_data; // @[SRAMTemplate.scala 76:26]
    end
    array_1__T_13_en_pipe_0 <= io_r_req_valid & _T;
    if (io_r_req_valid & _T) begin
      array_1__T_13_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if(array_2__T_9_en & array_2__T_9_mask) begin
      array_2[array_2__T_9_addr] <= array_2__T_9_data; // @[SRAMTemplate.scala 76:26]
    end
    array_2__T_13_en_pipe_0 <= io_r_req_valid & _T;
    if (io_r_req_valid & _T) begin
      array_2__T_13_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if(array_3__T_9_en & array_3__T_9_mask) begin
      array_3[array_3__T_9_addr] <= array_3__T_9_data; // @[SRAMTemplate.scala 76:26]
    end
    array_3__T_13_en_pipe_0 <= io_r_req_valid & _T;
    if (io_r_req_valid & _T) begin
      array_3__T_13_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
  end
endmodule
module Arbiter_3(
  output       io_in_0_ready,
  input        io_in_0_valid,
  input  [9:0] io_in_0_bits_setIdx,
  output       io_in_1_ready,
  input        io_in_1_valid,
  input  [9:0] io_in_1_bits_setIdx,
  input        io_out_ready,
  output       io_out_valid,
  output [9:0] io_out_bits_setIdx
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  wire  _T_2 = ~grant_1; // @[Arbiter.scala 135:19]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:14]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_out_valid = _T_2 | io_in_1_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
endmodule
module SRAMTemplateWithArbiter_1(
  input         clock,
  input         reset,
  output        io_r_0_req_ready,
  input         io_r_0_req_valid,
  input  [9:0]  io_r_0_req_bits_setIdx,
  output [63:0] io_r_0_resp_data_0_data,
  output [63:0] io_r_0_resp_data_1_data,
  output [63:0] io_r_0_resp_data_2_data,
  output [63:0] io_r_0_resp_data_3_data,
  output        io_r_1_req_ready,
  input         io_r_1_req_valid,
  input  [9:0]  io_r_1_req_bits_setIdx,
  output [63:0] io_r_1_resp_data_0_data,
  output [63:0] io_r_1_resp_data_1_data,
  output [63:0] io_r_1_resp_data_2_data,
  output [63:0] io_r_1_resp_data_3_data,
  input         io_w_req_valid,
  input  [9:0]  io_w_req_bits_setIdx,
  input  [63:0] io_w_req_bits_data_data,
  input  [3:0]  io_w_req_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  ram_clock; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_r_req_ready; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_r_req_valid; // @[SRAMTemplate.scala 121:19]
  wire [9:0] ram_io_r_req_bits_setIdx; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_r_resp_data_0_data; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_r_resp_data_1_data; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_r_resp_data_2_data; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_r_resp_data_3_data; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_w_req_valid; // @[SRAMTemplate.scala 121:19]
  wire [9:0] ram_io_w_req_bits_setIdx; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_w_req_bits_data_data; // @[SRAMTemplate.scala 121:19]
  wire [3:0] ram_io_w_req_bits_waymask; // @[SRAMTemplate.scala 121:19]
  wire  readArb_io_in_0_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_in_0_valid; // @[SRAMTemplate.scala 124:23]
  wire [9:0] readArb_io_in_0_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_in_1_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_in_1_valid; // @[SRAMTemplate.scala 124:23]
  wire [9:0] readArb_io_in_1_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_out_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_out_valid; // @[SRAMTemplate.scala 124:23]
  wire [9:0] readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  reg  _T_1; // @[SRAMTemplate.scala 130:58]
  reg [63:0] _T_3_0_data; // @[Reg.scala 27:20]
  reg [63:0] _T_3_1_data; // @[Reg.scala 27:20]
  reg [63:0] _T_3_2_data; // @[Reg.scala 27:20]
  reg [63:0] _T_3_3_data; // @[Reg.scala 27:20]
  reg  _T_6; // @[SRAMTemplate.scala 130:58]
  reg [63:0] _T_8_0_data; // @[Reg.scala 27:20]
  reg [63:0] _T_8_1_data; // @[Reg.scala 27:20]
  reg [63:0] _T_8_2_data; // @[Reg.scala 27:20]
  reg [63:0] _T_8_3_data; // @[Reg.scala 27:20]
  SRAMTemplate_2 ram ( // @[SRAMTemplate.scala 121:19]
    .clock(ram_clock),
    .io_r_req_ready(ram_io_r_req_ready),
    .io_r_req_valid(ram_io_r_req_valid),
    .io_r_req_bits_setIdx(ram_io_r_req_bits_setIdx),
    .io_r_resp_data_0_data(ram_io_r_resp_data_0_data),
    .io_r_resp_data_1_data(ram_io_r_resp_data_1_data),
    .io_r_resp_data_2_data(ram_io_r_resp_data_2_data),
    .io_r_resp_data_3_data(ram_io_r_resp_data_3_data),
    .io_w_req_valid(ram_io_w_req_valid),
    .io_w_req_bits_setIdx(ram_io_w_req_bits_setIdx),
    .io_w_req_bits_data_data(ram_io_w_req_bits_data_data),
    .io_w_req_bits_waymask(ram_io_w_req_bits_waymask)
  );
  Arbiter_3 readArb ( // @[SRAMTemplate.scala 124:23]
    .io_in_0_ready(readArb_io_in_0_ready),
    .io_in_0_valid(readArb_io_in_0_valid),
    .io_in_0_bits_setIdx(readArb_io_in_0_bits_setIdx),
    .io_in_1_ready(readArb_io_in_1_ready),
    .io_in_1_valid(readArb_io_in_1_valid),
    .io_in_1_bits_setIdx(readArb_io_in_1_bits_setIdx),
    .io_out_ready(readArb_io_out_ready),
    .io_out_valid(readArb_io_out_valid),
    .io_out_bits_setIdx(readArb_io_out_bits_setIdx)
  );
  assign io_r_0_req_ready = readArb_io_in_0_ready; // @[SRAMTemplate.scala 125:17]
  assign io_r_0_resp_data_0_data = _T_1 ? ram_io_r_resp_data_0_data : _T_3_0_data; // @[SRAMTemplate.scala 130:17]
  assign io_r_0_resp_data_1_data = _T_1 ? ram_io_r_resp_data_1_data : _T_3_1_data; // @[SRAMTemplate.scala 130:17]
  assign io_r_0_resp_data_2_data = _T_1 ? ram_io_r_resp_data_2_data : _T_3_2_data; // @[SRAMTemplate.scala 130:17]
  assign io_r_0_resp_data_3_data = _T_1 ? ram_io_r_resp_data_3_data : _T_3_3_data; // @[SRAMTemplate.scala 130:17]
  assign io_r_1_req_ready = readArb_io_in_1_ready; // @[SRAMTemplate.scala 125:17]
  assign io_r_1_resp_data_0_data = _T_6 ? ram_io_r_resp_data_0_data : _T_8_0_data; // @[SRAMTemplate.scala 130:17]
  assign io_r_1_resp_data_1_data = _T_6 ? ram_io_r_resp_data_1_data : _T_8_1_data; // @[SRAMTemplate.scala 130:17]
  assign io_r_1_resp_data_2_data = _T_6 ? ram_io_r_resp_data_2_data : _T_8_2_data; // @[SRAMTemplate.scala 130:17]
  assign io_r_1_resp_data_3_data = _T_6 ? ram_io_r_resp_data_3_data : _T_8_3_data; // @[SRAMTemplate.scala 130:17]
  assign ram_clock = clock;
  assign ram_io_r_req_valid = readArb_io_out_valid; // @[SRAMTemplate.scala 126:16]
  assign ram_io_r_req_bits_setIdx = readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 126:16]
  assign ram_io_w_req_valid = io_w_req_valid; // @[SRAMTemplate.scala 122:12]
  assign ram_io_w_req_bits_setIdx = io_w_req_bits_setIdx; // @[SRAMTemplate.scala 122:12]
  assign ram_io_w_req_bits_data_data = io_w_req_bits_data_data; // @[SRAMTemplate.scala 122:12]
  assign ram_io_w_req_bits_waymask = io_w_req_bits_waymask; // @[SRAMTemplate.scala 122:12]
  assign readArb_io_in_0_valid = io_r_0_req_valid; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_in_0_bits_setIdx = io_r_0_req_bits_setIdx; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_in_1_valid = io_r_1_req_valid; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_in_1_bits_setIdx = io_r_1_req_bits_setIdx; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_out_ready = ram_io_r_req_ready; // @[SRAMTemplate.scala 126:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1 = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  _T_3_0_data = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  _T_3_1_data = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  _T_3_2_data = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  _T_3_3_data = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  _T_6 = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  _T_8_0_data = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  _T_8_1_data = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  _T_8_2_data = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  _T_8_3_data = _RAND_9[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_1 <= io_r_0_req_ready & io_r_0_req_valid;
    if (reset) begin
      _T_3_0_data <= 64'h0;
    end else if (_T_1) begin
      _T_3_0_data <= ram_io_r_resp_data_0_data;
    end
    if (reset) begin
      _T_3_1_data <= 64'h0;
    end else if (_T_1) begin
      _T_3_1_data <= ram_io_r_resp_data_1_data;
    end
    if (reset) begin
      _T_3_2_data <= 64'h0;
    end else if (_T_1) begin
      _T_3_2_data <= ram_io_r_resp_data_2_data;
    end
    if (reset) begin
      _T_3_3_data <= 64'h0;
    end else if (_T_1) begin
      _T_3_3_data <= ram_io_r_resp_data_3_data;
    end
    _T_6 <= io_r_1_req_ready & io_r_1_req_valid;
    if (reset) begin
      _T_8_0_data <= 64'h0;
    end else if (_T_6) begin
      _T_8_0_data <= ram_io_r_resp_data_0_data;
    end
    if (reset) begin
      _T_8_1_data <= 64'h0;
    end else if (_T_6) begin
      _T_8_1_data <= ram_io_r_resp_data_1_data;
    end
    if (reset) begin
      _T_8_2_data <= 64'h0;
    end else if (_T_6) begin
      _T_8_2_data <= ram_io_r_resp_data_2_data;
    end
    if (reset) begin
      _T_8_3_data <= 64'h0;
    end else if (_T_6) begin
      _T_8_3_data <= ram_io_r_resp_data_3_data;
    end
  end
endmodule
module Arbiter_4(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input  [86:0] io_in_0_bits_user,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [86:0] io_out_bits_user
);
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:14]
  assign io_out_valid = io_in_0_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_addr = io_in_0_bits_addr; // @[Arbiter.scala 124:15]
  assign io_out_bits_user = io_in_0_bits_user; // @[Arbiter.scala 124:15]
endmodule
module Cache(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [86:0] io_in_req_bits_user,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  output [86:0] io_in_resp_bits_user,
  input  [1:0]  io_flush,
  input         io_out_mem_req_ready,
  output        io_out_mem_req_valid,
  output [31:0] io_out_mem_req_bits_addr,
  output [3:0]  io_out_mem_req_bits_cmd,
  output [63:0] io_out_mem_req_bits_wdata,
  input         io_out_mem_resp_valid,
  input  [3:0]  io_out_mem_resp_bits_cmd,
  input  [63:0] io_out_mem_resp_bits_rdata,
  input         io_mmio_req_ready,
  output        io_mmio_req_valid,
  output [31:0] io_mmio_req_bits_addr,
  input         io_mmio_resp_valid,
  input  [63:0] io_mmio_resp_bits_rdata,
  output        io_empty,
  input         MOUFlushICache,
  input         DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [95:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [95:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
`endif // RANDOMIZE_REG_INIT
  wire  s1_clock; // @[Cache.scala 475:18]
  wire  s1_reset; // @[Cache.scala 475:18]
  wire  s1_io_in_ready; // @[Cache.scala 475:18]
  wire  s1_io_in_valid; // @[Cache.scala 475:18]
  wire [31:0] s1_io_in_bits_addr; // @[Cache.scala 475:18]
  wire [2:0] s1_io_in_bits_size; // @[Cache.scala 475:18]
  wire [3:0] s1_io_in_bits_cmd; // @[Cache.scala 475:18]
  wire [7:0] s1_io_in_bits_wmask; // @[Cache.scala 475:18]
  wire [63:0] s1_io_in_bits_wdata; // @[Cache.scala 475:18]
  wire [86:0] s1_io_in_bits_user; // @[Cache.scala 475:18]
  wire  s1_io_out_ready; // @[Cache.scala 475:18]
  wire  s1_io_out_valid; // @[Cache.scala 475:18]
  wire [31:0] s1_io_out_bits_req_addr; // @[Cache.scala 475:18]
  wire [86:0] s1_io_out_bits_req_user; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_req_ready; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_req_valid; // @[Cache.scala 475:18]
  wire [6:0] s1_io_metaReadBus_req_bits_setIdx; // @[Cache.scala 475:18]
  wire [18:0] s1_io_metaReadBus_resp_data_0_tag; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_0_valid; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_0_dirty; // @[Cache.scala 475:18]
  wire [18:0] s1_io_metaReadBus_resp_data_1_tag; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_1_valid; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_1_dirty; // @[Cache.scala 475:18]
  wire [18:0] s1_io_metaReadBus_resp_data_2_tag; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_2_valid; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_2_dirty; // @[Cache.scala 475:18]
  wire [18:0] s1_io_metaReadBus_resp_data_3_tag; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_3_valid; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_3_dirty; // @[Cache.scala 475:18]
  wire  s1_io_dataReadBus_req_ready; // @[Cache.scala 475:18]
  wire  s1_io_dataReadBus_req_valid; // @[Cache.scala 475:18]
  wire [9:0] s1_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 475:18]
  wire [63:0] s1_io_dataReadBus_resp_data_0_data; // @[Cache.scala 475:18]
  wire [63:0] s1_io_dataReadBus_resp_data_1_data; // @[Cache.scala 475:18]
  wire [63:0] s1_io_dataReadBus_resp_data_2_data; // @[Cache.scala 475:18]
  wire [63:0] s1_io_dataReadBus_resp_data_3_data; // @[Cache.scala 475:18]
  wire  s1_DISPLAY_ENABLE; // @[Cache.scala 475:18]
  wire  s2_clock; // @[Cache.scala 476:18]
  wire  s2_reset; // @[Cache.scala 476:18]
  wire  s2_io_in_ready; // @[Cache.scala 476:18]
  wire  s2_io_in_valid; // @[Cache.scala 476:18]
  wire [31:0] s2_io_in_bits_req_addr; // @[Cache.scala 476:18]
  wire [2:0] s2_io_in_bits_req_size; // @[Cache.scala 476:18]
  wire [3:0] s2_io_in_bits_req_cmd; // @[Cache.scala 476:18]
  wire [7:0] s2_io_in_bits_req_wmask; // @[Cache.scala 476:18]
  wire [63:0] s2_io_in_bits_req_wdata; // @[Cache.scala 476:18]
  wire [86:0] s2_io_in_bits_req_user; // @[Cache.scala 476:18]
  wire  s2_io_out_ready; // @[Cache.scala 476:18]
  wire  s2_io_out_valid; // @[Cache.scala 476:18]
  wire [31:0] s2_io_out_bits_req_addr; // @[Cache.scala 476:18]
  wire [86:0] s2_io_out_bits_req_user; // @[Cache.scala 476:18]
  wire [18:0] s2_io_out_bits_metas_0_tag; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_0_valid; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_0_dirty; // @[Cache.scala 476:18]
  wire [18:0] s2_io_out_bits_metas_1_tag; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_1_valid; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_1_dirty; // @[Cache.scala 476:18]
  wire [18:0] s2_io_out_bits_metas_2_tag; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_2_valid; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_2_dirty; // @[Cache.scala 476:18]
  wire [18:0] s2_io_out_bits_metas_3_tag; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_3_valid; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_3_dirty; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_datas_0_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_datas_1_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_datas_2_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_datas_3_data; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_hit; // @[Cache.scala 476:18]
  wire [3:0] s2_io_out_bits_waymask; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_mmio; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_isForwardData; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_forwardData_data_data; // @[Cache.scala 476:18]
  wire [3:0] s2_io_out_bits_forwardData_waymask; // @[Cache.scala 476:18]
  wire [18:0] s2_io_metaReadResp_0_tag; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_0_valid; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_0_dirty; // @[Cache.scala 476:18]
  wire [18:0] s2_io_metaReadResp_1_tag; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_1_valid; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_1_dirty; // @[Cache.scala 476:18]
  wire [18:0] s2_io_metaReadResp_2_tag; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_2_valid; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_2_dirty; // @[Cache.scala 476:18]
  wire [18:0] s2_io_metaReadResp_3_tag; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_3_valid; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_3_dirty; // @[Cache.scala 476:18]
  wire [63:0] s2_io_dataReadResp_0_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_dataReadResp_1_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_dataReadResp_2_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_dataReadResp_3_data; // @[Cache.scala 476:18]
  wire  s2_io_metaWriteBus_req_valid; // @[Cache.scala 476:18]
  wire [6:0] s2_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 476:18]
  wire [18:0] s2_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 476:18]
  wire  s2_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 476:18]
  wire [3:0] s2_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 476:18]
  wire  s2_io_dataWriteBus_req_valid; // @[Cache.scala 476:18]
  wire [9:0] s2_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 476:18]
  wire [63:0] s2_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 476:18]
  wire [3:0] s2_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 476:18]
  wire  s2_DISPLAY_ENABLE; // @[Cache.scala 476:18]
  wire  s3_clock; // @[Cache.scala 477:18]
  wire  s3_reset; // @[Cache.scala 477:18]
  wire  s3_io_in_ready; // @[Cache.scala 477:18]
  wire  s3_io_in_valid; // @[Cache.scala 477:18]
  wire [31:0] s3_io_in_bits_req_addr; // @[Cache.scala 477:18]
  wire [2:0] s3_io_in_bits_req_size; // @[Cache.scala 477:18]
  wire [3:0] s3_io_in_bits_req_cmd; // @[Cache.scala 477:18]
  wire [7:0] s3_io_in_bits_req_wmask; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_req_wdata; // @[Cache.scala 477:18]
  wire [86:0] s3_io_in_bits_req_user; // @[Cache.scala 477:18]
  wire [18:0] s3_io_in_bits_metas_0_tag; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_0_valid; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_0_dirty; // @[Cache.scala 477:18]
  wire [18:0] s3_io_in_bits_metas_1_tag; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_1_valid; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_1_dirty; // @[Cache.scala 477:18]
  wire [18:0] s3_io_in_bits_metas_2_tag; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_2_valid; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_2_dirty; // @[Cache.scala 477:18]
  wire [18:0] s3_io_in_bits_metas_3_tag; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_3_valid; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_3_dirty; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_datas_0_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_datas_1_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_datas_2_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_datas_3_data; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_hit; // @[Cache.scala 477:18]
  wire [3:0] s3_io_in_bits_waymask; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_mmio; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_isForwardData; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_forwardData_data_data; // @[Cache.scala 477:18]
  wire [3:0] s3_io_in_bits_forwardData_waymask; // @[Cache.scala 477:18]
  wire  s3_io_out_ready; // @[Cache.scala 477:18]
  wire  s3_io_out_valid; // @[Cache.scala 477:18]
  wire [3:0] s3_io_out_bits_cmd; // @[Cache.scala 477:18]
  wire [63:0] s3_io_out_bits_rdata; // @[Cache.scala 477:18]
  wire [86:0] s3_io_out_bits_user; // @[Cache.scala 477:18]
  wire  s3_io_isFinish; // @[Cache.scala 477:18]
  wire  s3_io_flush; // @[Cache.scala 477:18]
  wire  s3_io_dataReadBus_req_ready; // @[Cache.scala 477:18]
  wire  s3_io_dataReadBus_req_valid; // @[Cache.scala 477:18]
  wire [9:0] s3_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 477:18]
  wire [63:0] s3_io_dataReadBus_resp_data_0_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_dataReadBus_resp_data_1_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_dataReadBus_resp_data_2_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_dataReadBus_resp_data_3_data; // @[Cache.scala 477:18]
  wire  s3_io_dataWriteBus_req_valid; // @[Cache.scala 477:18]
  wire [9:0] s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 477:18]
  wire [63:0] s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 477:18]
  wire [3:0] s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 477:18]
  wire  s3_io_metaWriteBus_req_valid; // @[Cache.scala 477:18]
  wire [6:0] s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 477:18]
  wire [18:0] s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 477:18]
  wire  s3_io_metaWriteBus_req_bits_data_valid; // @[Cache.scala 477:18]
  wire  s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 477:18]
  wire [3:0] s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 477:18]
  wire  s3_io_mem_req_ready; // @[Cache.scala 477:18]
  wire  s3_io_mem_req_valid; // @[Cache.scala 477:18]
  wire [31:0] s3_io_mem_req_bits_addr; // @[Cache.scala 477:18]
  wire [2:0] s3_io_mem_req_bits_size; // @[Cache.scala 477:18]
  wire [3:0] s3_io_mem_req_bits_cmd; // @[Cache.scala 477:18]
  wire [7:0] s3_io_mem_req_bits_wmask; // @[Cache.scala 477:18]
  wire [63:0] s3_io_mem_req_bits_wdata; // @[Cache.scala 477:18]
  wire  s3_io_mem_resp_ready; // @[Cache.scala 477:18]
  wire  s3_io_mem_resp_valid; // @[Cache.scala 477:18]
  wire [3:0] s3_io_mem_resp_bits_cmd; // @[Cache.scala 477:18]
  wire [63:0] s3_io_mem_resp_bits_rdata; // @[Cache.scala 477:18]
  wire  s3_io_mmio_req_ready; // @[Cache.scala 477:18]
  wire  s3_io_mmio_req_valid; // @[Cache.scala 477:18]
  wire [31:0] s3_io_mmio_req_bits_addr; // @[Cache.scala 477:18]
  wire  s3_io_mmio_resp_ready; // @[Cache.scala 477:18]
  wire  s3_io_mmio_resp_valid; // @[Cache.scala 477:18]
  wire [63:0] s3_io_mmio_resp_bits_rdata; // @[Cache.scala 477:18]
  wire  s3_io_cohResp_valid; // @[Cache.scala 477:18]
  wire  s3_DISPLAY_ENABLE; // @[Cache.scala 477:18]
  wire  metaArray_clock; // @[Cache.scala 478:25]
  wire  metaArray_reset; // @[Cache.scala 478:25]
  wire  metaArray_io_r_0_req_ready; // @[Cache.scala 478:25]
  wire  metaArray_io_r_0_req_valid; // @[Cache.scala 478:25]
  wire [6:0] metaArray_io_r_0_req_bits_setIdx; // @[Cache.scala 478:25]
  wire [18:0] metaArray_io_r_0_resp_data_0_tag; // @[Cache.scala 478:25]
  wire  metaArray_io_r_0_resp_data_0_valid; // @[Cache.scala 478:25]
  wire  metaArray_io_r_0_resp_data_0_dirty; // @[Cache.scala 478:25]
  wire [18:0] metaArray_io_r_0_resp_data_1_tag; // @[Cache.scala 478:25]
  wire  metaArray_io_r_0_resp_data_1_valid; // @[Cache.scala 478:25]
  wire  metaArray_io_r_0_resp_data_1_dirty; // @[Cache.scala 478:25]
  wire [18:0] metaArray_io_r_0_resp_data_2_tag; // @[Cache.scala 478:25]
  wire  metaArray_io_r_0_resp_data_2_valid; // @[Cache.scala 478:25]
  wire  metaArray_io_r_0_resp_data_2_dirty; // @[Cache.scala 478:25]
  wire [18:0] metaArray_io_r_0_resp_data_3_tag; // @[Cache.scala 478:25]
  wire  metaArray_io_r_0_resp_data_3_valid; // @[Cache.scala 478:25]
  wire  metaArray_io_r_0_resp_data_3_dirty; // @[Cache.scala 478:25]
  wire  metaArray_io_w_req_valid; // @[Cache.scala 478:25]
  wire [6:0] metaArray_io_w_req_bits_setIdx; // @[Cache.scala 478:25]
  wire [18:0] metaArray_io_w_req_bits_data_tag; // @[Cache.scala 478:25]
  wire  metaArray_io_w_req_bits_data_dirty; // @[Cache.scala 478:25]
  wire [3:0] metaArray_io_w_req_bits_waymask; // @[Cache.scala 478:25]
  wire  dataArray_clock; // @[Cache.scala 479:25]
  wire  dataArray_reset; // @[Cache.scala 479:25]
  wire  dataArray_io_r_0_req_ready; // @[Cache.scala 479:25]
  wire  dataArray_io_r_0_req_valid; // @[Cache.scala 479:25]
  wire [9:0] dataArray_io_r_0_req_bits_setIdx; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r_0_resp_data_0_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r_0_resp_data_1_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r_0_resp_data_2_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r_0_resp_data_3_data; // @[Cache.scala 479:25]
  wire  dataArray_io_r_1_req_ready; // @[Cache.scala 479:25]
  wire  dataArray_io_r_1_req_valid; // @[Cache.scala 479:25]
  wire [9:0] dataArray_io_r_1_req_bits_setIdx; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r_1_resp_data_0_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r_1_resp_data_1_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r_1_resp_data_2_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r_1_resp_data_3_data; // @[Cache.scala 479:25]
  wire  dataArray_io_w_req_valid; // @[Cache.scala 479:25]
  wire [9:0] dataArray_io_w_req_bits_setIdx; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_w_req_bits_data_data; // @[Cache.scala 479:25]
  wire [3:0] dataArray_io_w_req_bits_waymask; // @[Cache.scala 479:25]
  wire  arb_io_in_0_ready; // @[Cache.scala 488:19]
  wire  arb_io_in_0_valid; // @[Cache.scala 488:19]
  wire [31:0] arb_io_in_0_bits_addr; // @[Cache.scala 488:19]
  wire [86:0] arb_io_in_0_bits_user; // @[Cache.scala 488:19]
  wire  arb_io_out_ready; // @[Cache.scala 488:19]
  wire  arb_io_out_valid; // @[Cache.scala 488:19]
  wire [31:0] arb_io_out_bits_addr; // @[Cache.scala 488:19]
  wire [86:0] arb_io_out_bits_user; // @[Cache.scala 488:19]
  wire  _T_3 = s2_io_out_ready & s2_io_out_valid; // @[Decoupled.scala 40:37]
  reg  _T_5; // @[Pipeline.scala 24:24]
  wire  _GEN_0 = _T_3 ? 1'h0 : _T_5; // @[Pipeline.scala 25:25]
  wire  _T_6 = s1_io_out_valid & s2_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_1 = _T_6 | _GEN_0; // @[Pipeline.scala 26:38]
  reg [31:0] _T_8_req_addr; // @[Reg.scala 15:16]
  reg [86:0] _T_8_req_user; // @[Reg.scala 15:16]
  reg  _T_10; // @[Pipeline.scala 24:24]
  wire  _GEN_9 = s3_io_isFinish ? 1'h0 : _T_10; // @[Pipeline.scala 25:25]
  wire  _T_11 = s2_io_out_valid & s3_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_10 = _T_11 | _GEN_9; // @[Pipeline.scala 26:38]
  reg [31:0] _T_13_req_addr; // @[Reg.scala 15:16]
  reg [86:0] _T_13_req_user; // @[Reg.scala 15:16]
  reg [18:0] _T_13_metas_0_tag; // @[Reg.scala 15:16]
  reg  _T_13_metas_0_valid; // @[Reg.scala 15:16]
  reg  _T_13_metas_0_dirty; // @[Reg.scala 15:16]
  reg [18:0] _T_13_metas_1_tag; // @[Reg.scala 15:16]
  reg  _T_13_metas_1_valid; // @[Reg.scala 15:16]
  reg  _T_13_metas_1_dirty; // @[Reg.scala 15:16]
  reg [18:0] _T_13_metas_2_tag; // @[Reg.scala 15:16]
  reg  _T_13_metas_2_valid; // @[Reg.scala 15:16]
  reg  _T_13_metas_2_dirty; // @[Reg.scala 15:16]
  reg [18:0] _T_13_metas_3_tag; // @[Reg.scala 15:16]
  reg  _T_13_metas_3_valid; // @[Reg.scala 15:16]
  reg  _T_13_metas_3_dirty; // @[Reg.scala 15:16]
  reg [63:0] _T_13_datas_0_data; // @[Reg.scala 15:16]
  reg [63:0] _T_13_datas_1_data; // @[Reg.scala 15:16]
  reg [63:0] _T_13_datas_2_data; // @[Reg.scala 15:16]
  reg [63:0] _T_13_datas_3_data; // @[Reg.scala 15:16]
  reg  _T_13_hit; // @[Reg.scala 15:16]
  reg [3:0] _T_13_waymask; // @[Reg.scala 15:16]
  reg  _T_13_mmio; // @[Reg.scala 15:16]
  reg  _T_13_isForwardData; // @[Reg.scala 15:16]
  reg [63:0] _T_13_forwardData_data_data; // @[Reg.scala 15:16]
  reg [3:0] _T_13_forwardData_waymask; // @[Reg.scala 15:16]
  wire  _T_15 = ~s2_io_in_valid; // @[Cache.scala 503:15]
  wire  _T_16 = ~s3_io_in_valid; // @[Cache.scala 503:34]
  reg [63:0] _T_22; // @[GTimer.scala 24:20]
  wire [63:0] _T_24 = _T_22 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_28 = ~reset; // @[Debug.scala 56:24]
  reg [63:0] _T_31; // @[GTimer.scala 24:20]
  wire [63:0] _T_33 = _T_31 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_40; // @[GTimer.scala 24:20]
  wire [63:0] _T_42 = _T_40 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_49; // @[GTimer.scala 24:20]
  wire [63:0] _T_51 = _T_49 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_58; // @[GTimer.scala 24:20]
  wire [63:0] _T_60 = _T_58 + 64'h1; // @[GTimer.scala 25:12]
  wire  _GEN_41 = s1_io_in_valid & DISPLAY_ENABLE; // @[Debug.scala 56:24]
  wire  _GEN_43 = s2_io_in_valid & DISPLAY_ENABLE; // @[Debug.scala 56:24]
  wire  _GEN_45 = s3_io_in_valid & DISPLAY_ENABLE; // @[Debug.scala 56:24]
  CacheStage1 s1 ( // @[Cache.scala 475:18]
    .clock(s1_clock),
    .reset(s1_reset),
    .io_in_ready(s1_io_in_ready),
    .io_in_valid(s1_io_in_valid),
    .io_in_bits_addr(s1_io_in_bits_addr),
    .io_in_bits_size(s1_io_in_bits_size),
    .io_in_bits_cmd(s1_io_in_bits_cmd),
    .io_in_bits_wmask(s1_io_in_bits_wmask),
    .io_in_bits_wdata(s1_io_in_bits_wdata),
    .io_in_bits_user(s1_io_in_bits_user),
    .io_out_ready(s1_io_out_ready),
    .io_out_valid(s1_io_out_valid),
    .io_out_bits_req_addr(s1_io_out_bits_req_addr),
    .io_out_bits_req_user(s1_io_out_bits_req_user),
    .io_metaReadBus_req_ready(s1_io_metaReadBus_req_ready),
    .io_metaReadBus_req_valid(s1_io_metaReadBus_req_valid),
    .io_metaReadBus_req_bits_setIdx(s1_io_metaReadBus_req_bits_setIdx),
    .io_metaReadBus_resp_data_0_tag(s1_io_metaReadBus_resp_data_0_tag),
    .io_metaReadBus_resp_data_0_valid(s1_io_metaReadBus_resp_data_0_valid),
    .io_metaReadBus_resp_data_0_dirty(s1_io_metaReadBus_resp_data_0_dirty),
    .io_metaReadBus_resp_data_1_tag(s1_io_metaReadBus_resp_data_1_tag),
    .io_metaReadBus_resp_data_1_valid(s1_io_metaReadBus_resp_data_1_valid),
    .io_metaReadBus_resp_data_1_dirty(s1_io_metaReadBus_resp_data_1_dirty),
    .io_metaReadBus_resp_data_2_tag(s1_io_metaReadBus_resp_data_2_tag),
    .io_metaReadBus_resp_data_2_valid(s1_io_metaReadBus_resp_data_2_valid),
    .io_metaReadBus_resp_data_2_dirty(s1_io_metaReadBus_resp_data_2_dirty),
    .io_metaReadBus_resp_data_3_tag(s1_io_metaReadBus_resp_data_3_tag),
    .io_metaReadBus_resp_data_3_valid(s1_io_metaReadBus_resp_data_3_valid),
    .io_metaReadBus_resp_data_3_dirty(s1_io_metaReadBus_resp_data_3_dirty),
    .io_dataReadBus_req_ready(s1_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s1_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s1_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s1_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s1_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s1_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s1_io_dataReadBus_resp_data_3_data),
    .DISPLAY_ENABLE(s1_DISPLAY_ENABLE)
  );
  CacheStage2 s2 ( // @[Cache.scala 476:18]
    .clock(s2_clock),
    .reset(s2_reset),
    .io_in_ready(s2_io_in_ready),
    .io_in_valid(s2_io_in_valid),
    .io_in_bits_req_addr(s2_io_in_bits_req_addr),
    .io_in_bits_req_size(s2_io_in_bits_req_size),
    .io_in_bits_req_cmd(s2_io_in_bits_req_cmd),
    .io_in_bits_req_wmask(s2_io_in_bits_req_wmask),
    .io_in_bits_req_wdata(s2_io_in_bits_req_wdata),
    .io_in_bits_req_user(s2_io_in_bits_req_user),
    .io_out_ready(s2_io_out_ready),
    .io_out_valid(s2_io_out_valid),
    .io_out_bits_req_addr(s2_io_out_bits_req_addr),
    .io_out_bits_req_user(s2_io_out_bits_req_user),
    .io_out_bits_metas_0_tag(s2_io_out_bits_metas_0_tag),
    .io_out_bits_metas_0_valid(s2_io_out_bits_metas_0_valid),
    .io_out_bits_metas_0_dirty(s2_io_out_bits_metas_0_dirty),
    .io_out_bits_metas_1_tag(s2_io_out_bits_metas_1_tag),
    .io_out_bits_metas_1_valid(s2_io_out_bits_metas_1_valid),
    .io_out_bits_metas_1_dirty(s2_io_out_bits_metas_1_dirty),
    .io_out_bits_metas_2_tag(s2_io_out_bits_metas_2_tag),
    .io_out_bits_metas_2_valid(s2_io_out_bits_metas_2_valid),
    .io_out_bits_metas_2_dirty(s2_io_out_bits_metas_2_dirty),
    .io_out_bits_metas_3_tag(s2_io_out_bits_metas_3_tag),
    .io_out_bits_metas_3_valid(s2_io_out_bits_metas_3_valid),
    .io_out_bits_metas_3_dirty(s2_io_out_bits_metas_3_dirty),
    .io_out_bits_datas_0_data(s2_io_out_bits_datas_0_data),
    .io_out_bits_datas_1_data(s2_io_out_bits_datas_1_data),
    .io_out_bits_datas_2_data(s2_io_out_bits_datas_2_data),
    .io_out_bits_datas_3_data(s2_io_out_bits_datas_3_data),
    .io_out_bits_hit(s2_io_out_bits_hit),
    .io_out_bits_waymask(s2_io_out_bits_waymask),
    .io_out_bits_mmio(s2_io_out_bits_mmio),
    .io_out_bits_isForwardData(s2_io_out_bits_isForwardData),
    .io_out_bits_forwardData_data_data(s2_io_out_bits_forwardData_data_data),
    .io_out_bits_forwardData_waymask(s2_io_out_bits_forwardData_waymask),
    .io_metaReadResp_0_tag(s2_io_metaReadResp_0_tag),
    .io_metaReadResp_0_valid(s2_io_metaReadResp_0_valid),
    .io_metaReadResp_0_dirty(s2_io_metaReadResp_0_dirty),
    .io_metaReadResp_1_tag(s2_io_metaReadResp_1_tag),
    .io_metaReadResp_1_valid(s2_io_metaReadResp_1_valid),
    .io_metaReadResp_1_dirty(s2_io_metaReadResp_1_dirty),
    .io_metaReadResp_2_tag(s2_io_metaReadResp_2_tag),
    .io_metaReadResp_2_valid(s2_io_metaReadResp_2_valid),
    .io_metaReadResp_2_dirty(s2_io_metaReadResp_2_dirty),
    .io_metaReadResp_3_tag(s2_io_metaReadResp_3_tag),
    .io_metaReadResp_3_valid(s2_io_metaReadResp_3_valid),
    .io_metaReadResp_3_dirty(s2_io_metaReadResp_3_dirty),
    .io_dataReadResp_0_data(s2_io_dataReadResp_0_data),
    .io_dataReadResp_1_data(s2_io_dataReadResp_1_data),
    .io_dataReadResp_2_data(s2_io_dataReadResp_2_data),
    .io_dataReadResp_3_data(s2_io_dataReadResp_3_data),
    .io_metaWriteBus_req_valid(s2_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s2_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s2_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_data_dirty(s2_io_metaWriteBus_req_bits_data_dirty),
    .io_metaWriteBus_req_bits_waymask(s2_io_metaWriteBus_req_bits_waymask),
    .io_dataWriteBus_req_valid(s2_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s2_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s2_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s2_io_dataWriteBus_req_bits_waymask),
    .DISPLAY_ENABLE(s2_DISPLAY_ENABLE)
  );
  CacheStage3 s3 ( // @[Cache.scala 477:18]
    .clock(s3_clock),
    .reset(s3_reset),
    .io_in_ready(s3_io_in_ready),
    .io_in_valid(s3_io_in_valid),
    .io_in_bits_req_addr(s3_io_in_bits_req_addr),
    .io_in_bits_req_size(s3_io_in_bits_req_size),
    .io_in_bits_req_cmd(s3_io_in_bits_req_cmd),
    .io_in_bits_req_wmask(s3_io_in_bits_req_wmask),
    .io_in_bits_req_wdata(s3_io_in_bits_req_wdata),
    .io_in_bits_req_user(s3_io_in_bits_req_user),
    .io_in_bits_metas_0_tag(s3_io_in_bits_metas_0_tag),
    .io_in_bits_metas_0_valid(s3_io_in_bits_metas_0_valid),
    .io_in_bits_metas_0_dirty(s3_io_in_bits_metas_0_dirty),
    .io_in_bits_metas_1_tag(s3_io_in_bits_metas_1_tag),
    .io_in_bits_metas_1_valid(s3_io_in_bits_metas_1_valid),
    .io_in_bits_metas_1_dirty(s3_io_in_bits_metas_1_dirty),
    .io_in_bits_metas_2_tag(s3_io_in_bits_metas_2_tag),
    .io_in_bits_metas_2_valid(s3_io_in_bits_metas_2_valid),
    .io_in_bits_metas_2_dirty(s3_io_in_bits_metas_2_dirty),
    .io_in_bits_metas_3_tag(s3_io_in_bits_metas_3_tag),
    .io_in_bits_metas_3_valid(s3_io_in_bits_metas_3_valid),
    .io_in_bits_metas_3_dirty(s3_io_in_bits_metas_3_dirty),
    .io_in_bits_datas_0_data(s3_io_in_bits_datas_0_data),
    .io_in_bits_datas_1_data(s3_io_in_bits_datas_1_data),
    .io_in_bits_datas_2_data(s3_io_in_bits_datas_2_data),
    .io_in_bits_datas_3_data(s3_io_in_bits_datas_3_data),
    .io_in_bits_hit(s3_io_in_bits_hit),
    .io_in_bits_waymask(s3_io_in_bits_waymask),
    .io_in_bits_mmio(s3_io_in_bits_mmio),
    .io_in_bits_isForwardData(s3_io_in_bits_isForwardData),
    .io_in_bits_forwardData_data_data(s3_io_in_bits_forwardData_data_data),
    .io_in_bits_forwardData_waymask(s3_io_in_bits_forwardData_waymask),
    .io_out_ready(s3_io_out_ready),
    .io_out_valid(s3_io_out_valid),
    .io_out_bits_cmd(s3_io_out_bits_cmd),
    .io_out_bits_rdata(s3_io_out_bits_rdata),
    .io_out_bits_user(s3_io_out_bits_user),
    .io_isFinish(s3_io_isFinish),
    .io_flush(s3_io_flush),
    .io_dataReadBus_req_ready(s3_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s3_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s3_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s3_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s3_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s3_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s3_io_dataReadBus_resp_data_3_data),
    .io_dataWriteBus_req_valid(s3_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s3_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s3_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s3_io_dataWriteBus_req_bits_waymask),
    .io_metaWriteBus_req_valid(s3_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s3_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s3_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_data_valid(s3_io_metaWriteBus_req_bits_data_valid),
    .io_metaWriteBus_req_bits_data_dirty(s3_io_metaWriteBus_req_bits_data_dirty),
    .io_metaWriteBus_req_bits_waymask(s3_io_metaWriteBus_req_bits_waymask),
    .io_mem_req_ready(s3_io_mem_req_ready),
    .io_mem_req_valid(s3_io_mem_req_valid),
    .io_mem_req_bits_addr(s3_io_mem_req_bits_addr),
    .io_mem_req_bits_size(s3_io_mem_req_bits_size),
    .io_mem_req_bits_cmd(s3_io_mem_req_bits_cmd),
    .io_mem_req_bits_wmask(s3_io_mem_req_bits_wmask),
    .io_mem_req_bits_wdata(s3_io_mem_req_bits_wdata),
    .io_mem_resp_ready(s3_io_mem_resp_ready),
    .io_mem_resp_valid(s3_io_mem_resp_valid),
    .io_mem_resp_bits_cmd(s3_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_rdata(s3_io_mem_resp_bits_rdata),
    .io_mmio_req_ready(s3_io_mmio_req_ready),
    .io_mmio_req_valid(s3_io_mmio_req_valid),
    .io_mmio_req_bits_addr(s3_io_mmio_req_bits_addr),
    .io_mmio_resp_ready(s3_io_mmio_resp_ready),
    .io_mmio_resp_valid(s3_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(s3_io_mmio_resp_bits_rdata),
    .io_cohResp_valid(s3_io_cohResp_valid),
    .DISPLAY_ENABLE(s3_DISPLAY_ENABLE)
  );
  SRAMTemplateWithArbiter metaArray ( // @[Cache.scala 478:25]
    .clock(metaArray_clock),
    .reset(metaArray_reset),
    .io_r_0_req_ready(metaArray_io_r_0_req_ready),
    .io_r_0_req_valid(metaArray_io_r_0_req_valid),
    .io_r_0_req_bits_setIdx(metaArray_io_r_0_req_bits_setIdx),
    .io_r_0_resp_data_0_tag(metaArray_io_r_0_resp_data_0_tag),
    .io_r_0_resp_data_0_valid(metaArray_io_r_0_resp_data_0_valid),
    .io_r_0_resp_data_0_dirty(metaArray_io_r_0_resp_data_0_dirty),
    .io_r_0_resp_data_1_tag(metaArray_io_r_0_resp_data_1_tag),
    .io_r_0_resp_data_1_valid(metaArray_io_r_0_resp_data_1_valid),
    .io_r_0_resp_data_1_dirty(metaArray_io_r_0_resp_data_1_dirty),
    .io_r_0_resp_data_2_tag(metaArray_io_r_0_resp_data_2_tag),
    .io_r_0_resp_data_2_valid(metaArray_io_r_0_resp_data_2_valid),
    .io_r_0_resp_data_2_dirty(metaArray_io_r_0_resp_data_2_dirty),
    .io_r_0_resp_data_3_tag(metaArray_io_r_0_resp_data_3_tag),
    .io_r_0_resp_data_3_valid(metaArray_io_r_0_resp_data_3_valid),
    .io_r_0_resp_data_3_dirty(metaArray_io_r_0_resp_data_3_dirty),
    .io_w_req_valid(metaArray_io_w_req_valid),
    .io_w_req_bits_setIdx(metaArray_io_w_req_bits_setIdx),
    .io_w_req_bits_data_tag(metaArray_io_w_req_bits_data_tag),
    .io_w_req_bits_data_dirty(metaArray_io_w_req_bits_data_dirty),
    .io_w_req_bits_waymask(metaArray_io_w_req_bits_waymask)
  );
  SRAMTemplateWithArbiter_1 dataArray ( // @[Cache.scala 479:25]
    .clock(dataArray_clock),
    .reset(dataArray_reset),
    .io_r_0_req_ready(dataArray_io_r_0_req_ready),
    .io_r_0_req_valid(dataArray_io_r_0_req_valid),
    .io_r_0_req_bits_setIdx(dataArray_io_r_0_req_bits_setIdx),
    .io_r_0_resp_data_0_data(dataArray_io_r_0_resp_data_0_data),
    .io_r_0_resp_data_1_data(dataArray_io_r_0_resp_data_1_data),
    .io_r_0_resp_data_2_data(dataArray_io_r_0_resp_data_2_data),
    .io_r_0_resp_data_3_data(dataArray_io_r_0_resp_data_3_data),
    .io_r_1_req_ready(dataArray_io_r_1_req_ready),
    .io_r_1_req_valid(dataArray_io_r_1_req_valid),
    .io_r_1_req_bits_setIdx(dataArray_io_r_1_req_bits_setIdx),
    .io_r_1_resp_data_0_data(dataArray_io_r_1_resp_data_0_data),
    .io_r_1_resp_data_1_data(dataArray_io_r_1_resp_data_1_data),
    .io_r_1_resp_data_2_data(dataArray_io_r_1_resp_data_2_data),
    .io_r_1_resp_data_3_data(dataArray_io_r_1_resp_data_3_data),
    .io_w_req_valid(dataArray_io_w_req_valid),
    .io_w_req_bits_setIdx(dataArray_io_w_req_bits_setIdx),
    .io_w_req_bits_data_data(dataArray_io_w_req_bits_data_data),
    .io_w_req_bits_waymask(dataArray_io_w_req_bits_waymask)
  );
  Arbiter_4 arb ( // @[Cache.scala 488:19]
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_addr(arb_io_in_0_bits_addr),
    .io_in_0_bits_user(arb_io_in_0_bits_user),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_addr(arb_io_out_bits_addr),
    .io_out_bits_user(arb_io_out_bits_user)
  );
  assign io_in_req_ready = arb_io_in_0_ready; // @[Cache.scala 489:28]
  assign io_in_resp_valid = s3_io_out_valid; // @[Cache.scala 499:14 Cache.scala 505:20]
  assign io_in_resp_bits_rdata = s3_io_out_bits_rdata; // @[Cache.scala 499:14]
  assign io_in_resp_bits_user = s3_io_out_bits_user; // @[Cache.scala 499:14]
  assign io_out_mem_req_valid = s3_io_mem_req_valid; // @[Cache.scala 501:14]
  assign io_out_mem_req_bits_addr = s3_io_mem_req_bits_addr; // @[Cache.scala 501:14]
  assign io_out_mem_req_bits_cmd = s3_io_mem_req_bits_cmd; // @[Cache.scala 501:14]
  assign io_out_mem_req_bits_wdata = s3_io_mem_req_bits_wdata; // @[Cache.scala 501:14]
  assign io_mmio_req_valid = s3_io_mmio_req_valid; // @[Cache.scala 502:11]
  assign io_mmio_req_bits_addr = s3_io_mmio_req_bits_addr; // @[Cache.scala 502:11]
  assign io_empty = _T_15 & _T_16; // @[Cache.scala 503:12]
  assign s1_clock = clock;
  assign s1_reset = reset;
  assign s1_io_in_valid = arb_io_out_valid; // @[Cache.scala 491:12]
  assign s1_io_in_bits_addr = arb_io_out_bits_addr; // @[Cache.scala 491:12]
  assign s1_io_in_bits_size = 3'h3; // @[Cache.scala 491:12]
  assign s1_io_in_bits_cmd = 4'h0; // @[Cache.scala 491:12]
  assign s1_io_in_bits_wmask = 8'h0; // @[Cache.scala 491:12]
  assign s1_io_in_bits_wdata = 64'h0; // @[Cache.scala 491:12]
  assign s1_io_in_bits_user = arb_io_out_bits_user; // @[Cache.scala 491:12]
  assign s1_io_out_ready = s2_io_in_ready; // @[Pipeline.scala 29:16]
  assign s1_io_metaReadBus_req_ready = metaArray_io_r_0_req_ready; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_0_tag = metaArray_io_r_0_resp_data_0_tag; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_0_valid = metaArray_io_r_0_resp_data_0_valid; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_0_dirty = metaArray_io_r_0_resp_data_0_dirty; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_1_tag = metaArray_io_r_0_resp_data_1_tag; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_1_valid = metaArray_io_r_0_resp_data_1_valid; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_1_dirty = metaArray_io_r_0_resp_data_1_dirty; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_2_tag = metaArray_io_r_0_resp_data_2_tag; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_2_valid = metaArray_io_r_0_resp_data_2_valid; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_2_dirty = metaArray_io_r_0_resp_data_2_dirty; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_3_tag = metaArray_io_r_0_resp_data_3_tag; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_3_valid = metaArray_io_r_0_resp_data_3_valid; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_3_dirty = metaArray_io_r_0_resp_data_3_dirty; // @[Cache.scala 523:21]
  assign s1_io_dataReadBus_req_ready = dataArray_io_r_0_req_ready; // @[Cache.scala 524:21]
  assign s1_io_dataReadBus_resp_data_0_data = dataArray_io_r_0_resp_data_0_data; // @[Cache.scala 524:21]
  assign s1_io_dataReadBus_resp_data_1_data = dataArray_io_r_0_resp_data_1_data; // @[Cache.scala 524:21]
  assign s1_io_dataReadBus_resp_data_2_data = dataArray_io_r_0_resp_data_2_data; // @[Cache.scala 524:21]
  assign s1_io_dataReadBus_resp_data_3_data = dataArray_io_r_0_resp_data_3_data; // @[Cache.scala 524:21]
  assign s1_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign s2_clock = clock;
  assign s2_reset = reset;
  assign s2_io_in_valid = _T_5; // @[Pipeline.scala 31:17]
  assign s2_io_in_bits_req_addr = _T_8_req_addr; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_size = 3'h3; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_cmd = 4'h0; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_wmask = 8'h0; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_wdata = 64'h0; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_user = _T_8_req_user; // @[Pipeline.scala 30:16]
  assign s2_io_out_ready = s3_io_in_ready; // @[Pipeline.scala 29:16]
  assign s2_io_metaReadResp_0_tag = s1_io_metaReadBus_resp_data_0_tag; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_0_valid = s1_io_metaReadBus_resp_data_0_valid; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_0_dirty = s1_io_metaReadBus_resp_data_0_dirty; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_1_tag = s1_io_metaReadBus_resp_data_1_tag; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_1_valid = s1_io_metaReadBus_resp_data_1_valid; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_1_dirty = s1_io_metaReadBus_resp_data_1_dirty; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_2_tag = s1_io_metaReadBus_resp_data_2_tag; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_2_valid = s1_io_metaReadBus_resp_data_2_valid; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_2_dirty = s1_io_metaReadBus_resp_data_2_dirty; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_3_tag = s1_io_metaReadBus_resp_data_3_tag; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_3_valid = s1_io_metaReadBus_resp_data_3_valid; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_3_dirty = s1_io_metaReadBus_resp_data_3_dirty; // @[Cache.scala 530:22]
  assign s2_io_dataReadResp_0_data = s1_io_dataReadBus_resp_data_0_data; // @[Cache.scala 531:22]
  assign s2_io_dataReadResp_1_data = s1_io_dataReadBus_resp_data_1_data; // @[Cache.scala 531:22]
  assign s2_io_dataReadResp_2_data = s1_io_dataReadBus_resp_data_2_data; // @[Cache.scala 531:22]
  assign s2_io_dataReadResp_3_data = s1_io_dataReadBus_resp_data_3_data; // @[Cache.scala 531:22]
  assign s2_io_metaWriteBus_req_valid = s3_io_metaWriteBus_req_valid; // @[Cache.scala 533:22]
  assign s2_io_metaWriteBus_req_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 533:22]
  assign s2_io_metaWriteBus_req_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 533:22]
  assign s2_io_metaWriteBus_req_bits_data_dirty = s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 533:22]
  assign s2_io_metaWriteBus_req_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 533:22]
  assign s2_io_dataWriteBus_req_valid = s3_io_dataWriteBus_req_valid; // @[Cache.scala 532:22]
  assign s2_io_dataWriteBus_req_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 532:22]
  assign s2_io_dataWriteBus_req_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 532:22]
  assign s2_io_dataWriteBus_req_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 532:22]
  assign s2_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign s3_clock = clock;
  assign s3_reset = reset;
  assign s3_io_in_valid = _T_10; // @[Pipeline.scala 31:17]
  assign s3_io_in_bits_req_addr = _T_13_req_addr; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_size = 3'h3; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_cmd = 4'h0; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_wmask = 8'h0; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_wdata = 64'h0; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_user = _T_13_req_user; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_tag = _T_13_metas_0_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_valid = _T_13_metas_0_valid; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_dirty = _T_13_metas_0_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_tag = _T_13_metas_1_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_valid = _T_13_metas_1_valid; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_dirty = _T_13_metas_1_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_tag = _T_13_metas_2_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_valid = _T_13_metas_2_valid; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_dirty = _T_13_metas_2_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_tag = _T_13_metas_3_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_valid = _T_13_metas_3_valid; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_dirty = _T_13_metas_3_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_0_data = _T_13_datas_0_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_1_data = _T_13_datas_1_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_2_data = _T_13_datas_2_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_3_data = _T_13_datas_3_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_hit = _T_13_hit; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_waymask = _T_13_waymask; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_mmio = _T_13_mmio; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_isForwardData = _T_13_isForwardData; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_data_data = _T_13_forwardData_data_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_waymask = _T_13_forwardData_waymask; // @[Pipeline.scala 30:16]
  assign s3_io_out_ready = io_in_resp_ready; // @[Cache.scala 499:14]
  assign s3_io_flush = io_flush[1]; // @[Cache.scala 500:15]
  assign s3_io_dataReadBus_req_ready = dataArray_io_r_1_req_ready; // @[Cache.scala 525:21]
  assign s3_io_dataReadBus_resp_data_0_data = dataArray_io_r_1_resp_data_0_data; // @[Cache.scala 525:21]
  assign s3_io_dataReadBus_resp_data_1_data = dataArray_io_r_1_resp_data_1_data; // @[Cache.scala 525:21]
  assign s3_io_dataReadBus_resp_data_2_data = dataArray_io_r_1_resp_data_2_data; // @[Cache.scala 525:21]
  assign s3_io_dataReadBus_resp_data_3_data = dataArray_io_r_1_resp_data_3_data; // @[Cache.scala 525:21]
  assign s3_io_mem_req_ready = io_out_mem_req_ready; // @[Cache.scala 501:14]
  assign s3_io_mem_resp_valid = io_out_mem_resp_valid; // @[Cache.scala 501:14]
  assign s3_io_mem_resp_bits_cmd = io_out_mem_resp_bits_cmd; // @[Cache.scala 501:14]
  assign s3_io_mem_resp_bits_rdata = io_out_mem_resp_bits_rdata; // @[Cache.scala 501:14]
  assign s3_io_mmio_req_ready = io_mmio_req_ready; // @[Cache.scala 502:11]
  assign s3_io_mmio_resp_valid = io_mmio_resp_valid; // @[Cache.scala 502:11]
  assign s3_io_mmio_resp_bits_rdata = io_mmio_resp_bits_rdata; // @[Cache.scala 502:11]
  assign s3_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign metaArray_clock = clock;
  assign metaArray_reset = reset | MOUFlushICache; // @[Cache.scala 485:21]
  assign metaArray_io_r_0_req_valid = s1_io_metaReadBus_req_valid; // @[Cache.scala 523:21]
  assign metaArray_io_r_0_req_bits_setIdx = s1_io_metaReadBus_req_bits_setIdx; // @[Cache.scala 523:21]
  assign metaArray_io_w_req_valid = s3_io_metaWriteBus_req_valid; // @[Cache.scala 527:18]
  assign metaArray_io_w_req_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 527:18]
  assign metaArray_io_w_req_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 527:18]
  assign metaArray_io_w_req_bits_data_dirty = s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 527:18]
  assign metaArray_io_w_req_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 527:18]
  assign dataArray_clock = clock;
  assign dataArray_reset = reset;
  assign dataArray_io_r_0_req_valid = s1_io_dataReadBus_req_valid; // @[Cache.scala 524:21]
  assign dataArray_io_r_0_req_bits_setIdx = s1_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 524:21]
  assign dataArray_io_r_1_req_valid = s3_io_dataReadBus_req_valid; // @[Cache.scala 525:21]
  assign dataArray_io_r_1_req_bits_setIdx = s3_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 525:21]
  assign dataArray_io_w_req_valid = s3_io_dataWriteBus_req_valid; // @[Cache.scala 528:18]
  assign dataArray_io_w_req_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 528:18]
  assign dataArray_io_w_req_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 528:18]
  assign dataArray_io_w_req_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 528:18]
  assign arb_io_in_0_valid = io_in_req_valid; // @[Cache.scala 489:28]
  assign arb_io_in_0_bits_addr = io_in_req_bits_addr; // @[Cache.scala 489:28]
  assign arb_io_in_0_bits_user = io_in_req_bits_user; // @[Cache.scala 489:28]
  assign arb_io_out_ready = s1_io_in_ready; // @[Cache.scala 491:12]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_5 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _T_8_req_addr = _RAND_1[31:0];
  _RAND_2 = {3{`RANDOM}};
  _T_8_req_user = _RAND_2[86:0];
  _RAND_3 = {1{`RANDOM}};
  _T_10 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_13_req_addr = _RAND_4[31:0];
  _RAND_5 = {3{`RANDOM}};
  _T_13_req_user = _RAND_5[86:0];
  _RAND_6 = {1{`RANDOM}};
  _T_13_metas_0_tag = _RAND_6[18:0];
  _RAND_7 = {1{`RANDOM}};
  _T_13_metas_0_valid = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _T_13_metas_0_dirty = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _T_13_metas_1_tag = _RAND_9[18:0];
  _RAND_10 = {1{`RANDOM}};
  _T_13_metas_1_valid = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _T_13_metas_1_dirty = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _T_13_metas_2_tag = _RAND_12[18:0];
  _RAND_13 = {1{`RANDOM}};
  _T_13_metas_2_valid = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  _T_13_metas_2_dirty = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  _T_13_metas_3_tag = _RAND_15[18:0];
  _RAND_16 = {1{`RANDOM}};
  _T_13_metas_3_valid = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  _T_13_metas_3_dirty = _RAND_17[0:0];
  _RAND_18 = {2{`RANDOM}};
  _T_13_datas_0_data = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  _T_13_datas_1_data = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  _T_13_datas_2_data = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  _T_13_datas_3_data = _RAND_21[63:0];
  _RAND_22 = {1{`RANDOM}};
  _T_13_hit = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  _T_13_waymask = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  _T_13_mmio = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  _T_13_isForwardData = _RAND_25[0:0];
  _RAND_26 = {2{`RANDOM}};
  _T_13_forwardData_data_data = _RAND_26[63:0];
  _RAND_27 = {1{`RANDOM}};
  _T_13_forwardData_waymask = _RAND_27[3:0];
  _RAND_28 = {2{`RANDOM}};
  _T_22 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  _T_31 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  _T_40 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  _T_49 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  _T_58 = _RAND_32[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_5 <= 1'h0;
    end else if (io_flush[0]) begin
      _T_5 <= 1'h0;
    end else begin
      _T_5 <= _GEN_1;
    end
    if (_T_6) begin
      _T_8_req_addr <= s1_io_out_bits_req_addr;
    end
    if (_T_6) begin
      _T_8_req_user <= s1_io_out_bits_req_user;
    end
    if (reset) begin
      _T_10 <= 1'h0;
    end else if (io_flush[1]) begin
      _T_10 <= 1'h0;
    end else begin
      _T_10 <= _GEN_10;
    end
    if (_T_11) begin
      _T_13_req_addr <= s2_io_out_bits_req_addr;
    end
    if (_T_11) begin
      _T_13_req_user <= s2_io_out_bits_req_user;
    end
    if (_T_11) begin
      _T_13_metas_0_tag <= s2_io_out_bits_metas_0_tag;
    end
    if (_T_11) begin
      _T_13_metas_0_valid <= s2_io_out_bits_metas_0_valid;
    end
    if (_T_11) begin
      _T_13_metas_0_dirty <= s2_io_out_bits_metas_0_dirty;
    end
    if (_T_11) begin
      _T_13_metas_1_tag <= s2_io_out_bits_metas_1_tag;
    end
    if (_T_11) begin
      _T_13_metas_1_valid <= s2_io_out_bits_metas_1_valid;
    end
    if (_T_11) begin
      _T_13_metas_1_dirty <= s2_io_out_bits_metas_1_dirty;
    end
    if (_T_11) begin
      _T_13_metas_2_tag <= s2_io_out_bits_metas_2_tag;
    end
    if (_T_11) begin
      _T_13_metas_2_valid <= s2_io_out_bits_metas_2_valid;
    end
    if (_T_11) begin
      _T_13_metas_2_dirty <= s2_io_out_bits_metas_2_dirty;
    end
    if (_T_11) begin
      _T_13_metas_3_tag <= s2_io_out_bits_metas_3_tag;
    end
    if (_T_11) begin
      _T_13_metas_3_valid <= s2_io_out_bits_metas_3_valid;
    end
    if (_T_11) begin
      _T_13_metas_3_dirty <= s2_io_out_bits_metas_3_dirty;
    end
    if (_T_11) begin
      _T_13_datas_0_data <= s2_io_out_bits_datas_0_data;
    end
    if (_T_11) begin
      _T_13_datas_1_data <= s2_io_out_bits_datas_1_data;
    end
    if (_T_11) begin
      _T_13_datas_2_data <= s2_io_out_bits_datas_2_data;
    end
    if (_T_11) begin
      _T_13_datas_3_data <= s2_io_out_bits_datas_3_data;
    end
    if (_T_11) begin
      _T_13_hit <= s2_io_out_bits_hit;
    end
    if (_T_11) begin
      _T_13_waymask <= s2_io_out_bits_waymask;
    end
    if (_T_11) begin
      _T_13_mmio <= s2_io_out_bits_mmio;
    end
    if (_T_11) begin
      _T_13_isForwardData <= s2_io_out_bits_isForwardData;
    end
    if (_T_11) begin
      _T_13_forwardData_data_data <= s2_io_out_bits_forwardData_data_data;
    end
    if (_T_11) begin
      _T_13_forwardData_waymask <= s2_io_out_bits_forwardData_waymask;
    end
    if (reset) begin
      _T_22 <= 64'h0;
    end else begin
      _T_22 <= _T_24;
    end
    if (reset) begin
      _T_31 <= 64'h0;
    end else begin
      _T_31 <= _T_33;
    end
    if (reset) begin
      _T_40 <= 64'h0;
    end else begin
      _T_40 <= _T_42;
    end
    if (reset) begin
      _T_49 <= 64'h0;
    end else begin
      _T_49 <= _T_51;
    end
    if (reset) begin
      _T_58 <= 64'h0;
    end else begin
      _T_58 <= _T_60;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_28) begin
          $fwrite(32'h80000002,"[%d] Cache: ",_T_22); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_28) begin
          $fwrite(32'h80000002,"InReq(%d, %d) InResp(%d, %d) \n",io_in_req_valid,io_in_req_ready,io_in_resp_valid,io_in_resp_ready); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_28) begin
          $fwrite(32'h80000002,"[%d] Cache: ",_T_31); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_28) begin
          $fwrite(32'h80000002,"{IN s1:(%d,%d), s2:(%d,%d), s3:(%d,%d)} {OUT s1:(%d,%d), s2:(%d,%d), s3:(%d,%d)}\n",s1_io_in_valid,s1_io_in_ready,s2_io_in_valid,s2_io_in_ready,s3_io_in_valid,s3_io_in_ready,s1_io_out_valid,s1_io_out_ready,s2_io_out_valid,s2_io_out_ready,s3_io_out_valid,s3_io_out_ready); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_28) begin
          $fwrite(32'h80000002,"[%d] Cache: ",_T_40); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_28) begin
          $fwrite(32'h80000002,"[icache.S1]: addr = 0x%x, cmd = %d, size = %d, wmask = 0x%x, wdata = 0x%x\n",s1_io_in_bits_addr,s1_io_in_bits_cmd,s1_io_in_bits_size,s1_io_in_bits_wmask,s1_io_in_bits_wdata); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_43 & _T_28) begin
          $fwrite(32'h80000002,"[%d] Cache: ",_T_49); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_43 & _T_28) begin
          $fwrite(32'h80000002,"[icache.S2]: addr = 0x%x, cmd = %d, size = %d, wmask = 0x%x, wdata = 0x%x\n",s2_io_in_bits_req_addr,s2_io_in_bits_req_cmd,s2_io_in_bits_req_size,s2_io_in_bits_req_wmask,s2_io_in_bits_req_wdata); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_45 & _T_28) begin
          $fwrite(32'h80000002,"[%d] Cache: ",_T_58); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_45 & _T_28) begin
          $fwrite(32'h80000002,"[icache.S3]: addr = 0x%x, cmd = %d, size = %d, wmask = 0x%x, wdata = 0x%x\n",s3_io_in_bits_req_addr,s3_io_in_bits_req_cmd,s3_io_in_bits_req_size,s3_io_in_bits_req_wmask,s3_io_in_bits_req_wdata); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module EmbeddedTLBExec_1(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [38:0]  io_in_bits_addr,
  input  [2:0]   io_in_bits_size,
  input  [3:0]   io_in_bits_cmd,
  input  [7:0]   io_in_bits_wmask,
  input  [63:0]  io_in_bits_wdata,
  input          io_out_ready,
  output         io_out_valid,
  output [31:0]  io_out_bits_addr,
  output [2:0]   io_out_bits_size,
  output [3:0]   io_out_bits_cmd,
  output [7:0]   io_out_bits_wmask,
  output [63:0]  io_out_bits_wdata,
  input  [120:0] io_md_0,
  input  [120:0] io_md_1,
  input  [120:0] io_md_2,
  input  [120:0] io_md_3,
  output         io_mdWrite_wen,
  output [3:0]   io_mdWrite_windex,
  output [3:0]   io_mdWrite_waymask,
  output [120:0] io_mdWrite_wdata,
  input          io_mdReady,
  input          io_mem_req_ready,
  output         io_mem_req_valid,
  output [31:0]  io_mem_req_bits_addr,
  output [2:0]   io_mem_req_bits_size,
  output [3:0]   io_mem_req_bits_cmd,
  output [7:0]   io_mem_req_bits_wmask,
  output [63:0]  io_mem_req_bits_wdata,
  output         io_mem_resp_ready,
  input          io_mem_resp_valid,
  input  [3:0]   io_mem_resp_bits_cmd,
  input  [63:0]  io_mem_resp_bits_rdata,
  input  [63:0]  io_satp,
  input  [1:0]   io_pf_priviledgeMode,
  input          io_pf_status_sum,
  input          io_pf_status_mxr,
  output         io_pf_loadPF,
  output         io_pf_storePF,
  output [38:0]  io_pf_addr,
  output         io_ipf,
  output         io_isFinish,
  input          ISAMO,
  input          DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
`endif // RANDOMIZE_REG_INIT
  wire [8:0] vpn_vpn0 = io_in_bits_addr[20:12]; // @[EmbeddedTLB.scala 193:54]
  wire [8:0] vpn_vpn1 = io_in_bits_addr[29:21]; // @[EmbeddedTLB.scala 193:54]
  wire [8:0] vpn_vpn2 = io_in_bits_addr[38:30]; // @[EmbeddedTLB.scala 193:54]
  wire [19:0] satp_ppn = io_satp[19:0]; // @[EmbeddedTLB.scala 195:30]
  wire [15:0] satp_asid = io_satp[59:44]; // @[EmbeddedTLB.scala 195:30]
  wire  _T_39 = io_md_0[93:78] == satp_asid; // @[EmbeddedTLB.scala 204:117]
  wire  _T_40 = io_md_0[52] & _T_39; // @[EmbeddedTLB.scala 204:86]
  wire [17:0] _T_57 = {vpn_vpn2,vpn_vpn1}; // @[EmbeddedTLB.scala 204:201]
  wire [26:0] _T_58 = {vpn_vpn2,vpn_vpn1,vpn_vpn0}; // @[EmbeddedTLB.scala 204:201]
  wire [26:0] _T_59 = {9'h1ff,io_md_0[77:60]}; // @[Cat.scala 29:58]
  wire [26:0] _T_60 = _T_59 & io_md_0[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_62 = _T_59 & _T_58; // @[TLB.scala 131:84]
  wire  _T_63 = _T_60 == _T_62; // @[TLB.scala 131:48]
  wire  _T_64 = _T_40 & _T_63; // @[EmbeddedTLB.scala 204:132]
  wire  _T_91 = io_md_1[93:78] == satp_asid; // @[EmbeddedTLB.scala 204:117]
  wire  _T_92 = io_md_1[52] & _T_91; // @[EmbeddedTLB.scala 204:86]
  wire [26:0] _T_111 = {9'h1ff,io_md_1[77:60]}; // @[Cat.scala 29:58]
  wire [26:0] _T_112 = _T_111 & io_md_1[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_114 = _T_111 & _T_58; // @[TLB.scala 131:84]
  wire  _T_115 = _T_112 == _T_114; // @[TLB.scala 131:48]
  wire  _T_116 = _T_92 & _T_115; // @[EmbeddedTLB.scala 204:132]
  wire  _T_143 = io_md_2[93:78] == satp_asid; // @[EmbeddedTLB.scala 204:117]
  wire  _T_144 = io_md_2[52] & _T_143; // @[EmbeddedTLB.scala 204:86]
  wire [26:0] _T_163 = {9'h1ff,io_md_2[77:60]}; // @[Cat.scala 29:58]
  wire [26:0] _T_164 = _T_163 & io_md_2[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_166 = _T_163 & _T_58; // @[TLB.scala 131:84]
  wire  _T_167 = _T_164 == _T_166; // @[TLB.scala 131:48]
  wire  _T_168 = _T_144 & _T_167; // @[EmbeddedTLB.scala 204:132]
  wire  _T_195 = io_md_3[93:78] == satp_asid; // @[EmbeddedTLB.scala 204:117]
  wire  _T_196 = io_md_3[52] & _T_195; // @[EmbeddedTLB.scala 204:86]
  wire [26:0] _T_215 = {9'h1ff,io_md_3[77:60]}; // @[Cat.scala 29:58]
  wire [26:0] _T_216 = _T_215 & io_md_3[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_218 = _T_215 & _T_58; // @[TLB.scala 131:84]
  wire  _T_219 = _T_216 == _T_218; // @[TLB.scala 131:48]
  wire  _T_220 = _T_196 & _T_219; // @[EmbeddedTLB.scala 204:132]
  wire [3:0] hitVec = {_T_220,_T_168,_T_116,_T_64}; // @[EmbeddedTLB.scala 204:211]
  wire  _T_224 = |hitVec; // @[EmbeddedTLB.scala 205:35]
  wire  hit = io_in_valid & _T_224; // @[EmbeddedTLB.scala 205:25]
  wire  _T_226 = ~_T_224; // @[EmbeddedTLB.scala 206:29]
  wire  miss = io_in_valid & _T_226; // @[EmbeddedTLB.scala 206:26]
  reg [63:0] _T_227; // @[LFSR64.scala 25:23]
  wire  _T_230 = _T_227[0] ^ _T_227[1]; // @[LFSR64.scala 26:23]
  wire  _T_232 = _T_230 ^ _T_227[3]; // @[LFSR64.scala 26:33]
  wire  _T_234 = _T_232 ^ _T_227[4]; // @[LFSR64.scala 26:43]
  wire  _T_235 = _T_227 == 64'h0; // @[LFSR64.scala 28:24]
  wire [63:0] _T_237 = {_T_234,_T_227[63:1]}; // @[Cat.scala 29:58]
  wire [3:0] victimWaymask = 4'h1 << _T_227[1:0]; // @[EmbeddedTLB.scala 208:42]
  wire [3:0] waymask = hit ? hitVec : victimWaymask; // @[EmbeddedTLB.scala 209:20]
  wire [120:0] _T_244 = waymask[0] ? io_md_0 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_245 = waymask[1] ? io_md_1 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_246 = waymask[2] ? io_md_2 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_247 = waymask[3] ? io_md_3 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_248 = _T_244 | _T_245; // @[Mux.scala 27:72]
  wire [120:0] _T_249 = _T_248 | _T_246; // @[Mux.scala 27:72]
  wire [120:0] _T_250 = _T_249 | _T_247; // @[Mux.scala 27:72]
  wire [7:0] hitMeta_flag = _T_250[59:52]; // @[EmbeddedTLB.scala 215:70]
  wire [17:0] hitMeta_mask = _T_250[77:60]; // @[EmbeddedTLB.scala 215:70]
  wire [15:0] hitMeta_asid = _T_250[93:78]; // @[EmbeddedTLB.scala 215:70]
  wire [26:0] hitMeta_vpn = _T_250[120:94]; // @[EmbeddedTLB.scala 215:70]
  wire [31:0] hitData_pteaddr = _T_250[31:0]; // @[EmbeddedTLB.scala 216:70]
  wire [19:0] hitData_ppn = _T_250[51:32]; // @[EmbeddedTLB.scala 216:70]
  wire  hitFlag_v = hitMeta_flag[0]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_r = hitMeta_flag[1]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_w = hitMeta_flag[2]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_x = hitMeta_flag[3]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_u = hitMeta_flag[4]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_g = hitMeta_flag[5]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_a = hitMeta_flag[6]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_d = hitMeta_flag[7]; // @[EmbeddedTLB.scala 217:38]
  wire  _T_289 = ~hitFlag_a; // @[EmbeddedTLB.scala 221:23]
  wire  _T_290 = ~hitFlag_d; // @[EmbeddedTLB.scala 221:37]
  wire  _T_292 = _T_290 & io_in_bits_cmd[0]; // @[EmbeddedTLB.scala 221:48]
  wire  _T_293 = _T_289 | _T_292; // @[EmbeddedTLB.scala 221:34]
  wire  _T_294 = hit & _T_293; // @[EmbeddedTLB.scala 221:19]
  reg [2:0] state; // @[EmbeddedTLB.scala 247:22]
  wire  _T_370 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_314 = io_pf_priviledgeMode == 2'h0; // @[EmbeddedTLB.scala 226:62]
  wire  _T_315 = ~hitFlag_u; // @[EmbeddedTLB.scala 226:75]
  wire  _T_316 = _T_314 & _T_315; // @[EmbeddedTLB.scala 226:72]
  wire  _T_317 = ~_T_316; // @[EmbeddedTLB.scala 226:42]
  wire  _T_318 = hit & _T_317; // @[EmbeddedTLB.scala 226:39]
  wire  _T_319 = io_pf_priviledgeMode == 2'h1; // @[EmbeddedTLB.scala 226:110]
  wire  _T_320 = _T_319 & hitFlag_u; // @[EmbeddedTLB.scala 226:120]
  wire  _T_321 = ~io_pf_status_sum; // @[EmbeddedTLB.scala 226:137]
  wire  _T_323 = _T_320 & _T_321; // @[EmbeddedTLB.scala 226:133]
  wire  _T_324 = ~_T_323; // @[EmbeddedTLB.scala 226:90]
  wire  hitCheck = _T_318 & _T_324; // @[EmbeddedTLB.scala 226:87]
  wire  _T_325 = io_pf_status_mxr & hitFlag_x; // @[EmbeddedTLB.scala 228:57]
  wire  _T_326 = hitFlag_r | _T_325; // @[EmbeddedTLB.scala 228:40]
  wire  hitLoad = hitCheck & _T_326; // @[EmbeddedTLB.scala 228:26]
  wire  _T_329 = ~hitLoad; // @[EmbeddedTLB.scala 241:15]
  wire  _T_331 = ~io_in_bits_cmd[0]; // @[SimpleBus.scala 73:18]
  wire  _T_333 = ~io_in_bits_cmd[3]; // @[SimpleBus.scala 73:29]
  wire  _T_334 = _T_331 & _T_333; // @[SimpleBus.scala 73:26]
  wire  _T_335 = _T_329 & _T_334; // @[EmbeddedTLB.scala 241:24]
  wire  _T_336 = _T_335 & hit; // @[EmbeddedTLB.scala 241:40]
  wire  _T_337 = ~ISAMO; // @[EmbeddedTLB.scala 241:50]
  wire  _T_338 = _T_336 & _T_337; // @[EmbeddedTLB.scala 241:47]
  wire  _T_377 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_379 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_397 = io_mem_resp_ready & io_mem_resp_valid; // @[Decoupled.scala 40:37]
  wire  memRdata_flag_d = io_mem_resp_bits_rdata[7]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_a = io_mem_resp_bits_rdata[6]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_g = io_mem_resp_bits_rdata[5]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_u = io_mem_resp_bits_rdata[4]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_x = io_mem_resp_bits_rdata[3]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_w = io_mem_resp_bits_rdata[2]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_r = io_mem_resp_bits_rdata[1]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_v = io_mem_resp_bits_rdata[0]; // @[EmbeddedTLB.scala 255:49]
  wire [7:0] _T_387 = {memRdata_flag_d,memRdata_flag_a,memRdata_flag_g,memRdata_flag_u,memRdata_flag_x,memRdata_flag_w,memRdata_flag_r,memRdata_flag_v}; // @[EmbeddedTLB.scala 292:44]
  wire  _T_398 = _T_387[1] | _T_387[3]; // @[EmbeddedTLB.scala 297:34]
  wire  _T_399 = ~_T_398; // @[EmbeddedTLB.scala 297:21]
  reg [1:0] level; // @[EmbeddedTLB.scala 248:22]
  wire  _T_400 = level == 2'h3; // @[EmbeddedTLB.scala 297:58]
  wire  _T_401 = level == 2'h2; // @[EmbeddedTLB.scala 297:73]
  wire  _T_402 = _T_400 | _T_401; // @[EmbeddedTLB.scala 297:65]
  wire  _T_403 = _T_399 & _T_402; // @[EmbeddedTLB.scala 297:49]
  wire  _T_404 = ~_T_387[0]; // @[EmbeddedTLB.scala 298:16]
  wire  _T_405 = ~_T_387[1]; // @[EmbeddedTLB.scala 298:32]
  wire  _T_406 = _T_405 & _T_387[2]; // @[EmbeddedTLB.scala 298:44]
  wire  _T_407 = _T_404 | _T_406; // @[EmbeddedTLB.scala 298:28]
  wire  _T_414 = _T_334 & _T_337; // @[EmbeddedTLB.scala 302:38]
  wire  _GEN_19 = _T_407 ? _T_414 : _T_338; // @[EmbeddedTLB.scala 298:60]
  wire  _T_451 = level != 2'h0; // @[EmbeddedTLB.scala 313:27]
  wire  _T_453 = ~_T_387[4]; // @[EmbeddedTLB.scala 314:74]
  wire  _T_454 = _T_314 & _T_453; // @[EmbeddedTLB.scala 314:71]
  wire  _T_455 = ~_T_454; // @[EmbeddedTLB.scala 314:41]
  wire  _T_456 = _T_387[0] & _T_455; // @[EmbeddedTLB.scala 314:38]
  wire  _T_458 = _T_319 & _T_387[4]; // @[EmbeddedTLB.scala 314:120]
  wire  _T_461 = _T_458 & _T_321; // @[EmbeddedTLB.scala 314:134]
  wire  _T_462 = ~_T_461; // @[EmbeddedTLB.scala 314:90]
  wire  _T_463 = _T_456 & _T_462; // @[EmbeddedTLB.scala 314:87]
  wire  _T_465 = io_pf_status_mxr & _T_387[3]; // @[EmbeddedTLB.scala 316:68]
  wire  _T_466 = _T_387[1] | _T_465; // @[EmbeddedTLB.scala 316:51]
  wire  _T_467 = _T_463 & _T_466; // @[EmbeddedTLB.scala 316:36]
  wire  _T_485 = ~_T_467; // @[EmbeddedTLB.scala 330:19]
  wire  _T_491 = _T_485 & _T_334; // @[EmbeddedTLB.scala 330:29]
  wire  _T_468 = _T_463 & _T_387[2]; // @[EmbeddedTLB.scala 317:37]
  wire  _T_492 = ~_T_468; // @[EmbeddedTLB.scala 330:50]
  wire  _T_494 = _T_492 & io_in_bits_cmd[0]; // @[EmbeddedTLB.scala 330:61]
  wire  _T_495 = _T_491 | _T_494; // @[EmbeddedTLB.scala 330:46]
  wire  _GEN_23 = _T_495 ? _T_414 : _T_338; // @[EmbeddedTLB.scala 330:80]
  wire  _GEN_29 = _T_451 ? _GEN_23 : _T_338; // @[EmbeddedTLB.scala 313:36]
  wire  _GEN_35 = _T_403 ? _GEN_19 : _GEN_29; // @[EmbeddedTLB.scala 297:82]
  wire  _GEN_54 = _T_397 ? _GEN_35 : _T_338; // @[EmbeddedTLB.scala 293:33]
  wire  _GEN_78 = _T_379 ? _GEN_54 : _T_338; // @[Conditional.scala 39:67]
  wire  _GEN_91 = _T_377 ? _T_338 : _GEN_78; // @[Conditional.scala 39:67]
  wire  loadPF = _T_370 ? _T_338 : _GEN_91; // @[Conditional.scala 40:58]
  wire  hitStore = hitCheck & hitFlag_w; // @[EmbeddedTLB.scala 229:27]
  wire  _T_339 = ~hitStore; // @[EmbeddedTLB.scala 242:17]
  wire  _T_341 = _T_339 & io_in_bits_cmd[0]; // @[EmbeddedTLB.scala 242:27]
  wire  _T_342 = _T_341 & hit; // @[EmbeddedTLB.scala 242:44]
  wire  _T_351 = _T_336 & ISAMO; // @[EmbeddedTLB.scala 242:88]
  wire  _T_352 = _T_342 | _T_351; // @[EmbeddedTLB.scala 242:52]
  wire  _T_416 = io_in_bits_cmd[0] | ISAMO; // @[EmbeddedTLB.scala 303:40]
  wire  _GEN_20 = _T_407 ? _T_416 : _T_352; // @[EmbeddedTLB.scala 298:60]
  wire  _GEN_24 = _T_495 ? _T_416 : _T_352; // @[EmbeddedTLB.scala 330:80]
  wire  _GEN_30 = _T_451 ? _GEN_24 : _T_352; // @[EmbeddedTLB.scala 313:36]
  wire  _GEN_36 = _T_403 ? _GEN_20 : _GEN_30; // @[EmbeddedTLB.scala 297:82]
  wire  _GEN_55 = _T_397 ? _GEN_36 : _T_352; // @[EmbeddedTLB.scala 293:33]
  wire  _GEN_79 = _T_379 ? _GEN_55 : _T_352; // @[Conditional.scala 39:67]
  wire  _GEN_92 = _T_377 ? _T_352 : _GEN_79; // @[Conditional.scala 39:67]
  wire  storePF = _T_370 ? _T_352 : _GEN_92; // @[Conditional.scala 40:58]
  wire  _T_297 = loadPF | storePF; // @[EmbeddedTLB.scala 221:93]
  wire  _T_298 = io_pf_loadPF | io_pf_storePF; // @[Bundle.scala 135:23]
  wire  _T_299 = _T_297 | _T_298; // @[EmbeddedTLB.scala 221:104]
  wire  _T_300 = ~_T_299; // @[EmbeddedTLB.scala 221:84]
  wire  hitWB = _T_294 & _T_300; // @[EmbeddedTLB.scala 221:81]
  wire [7:0] _T_303 = {io_in_bits_cmd[0],1'h1,6'h0}; // @[Cat.scala 29:58]
  wire [7:0] _T_310 = {hitFlag_d,hitFlag_a,hitFlag_g,hitFlag_u,hitFlag_x,hitFlag_w,hitFlag_r,hitFlag_v}; // @[EmbeddedTLB.scala 222:79]
  wire [7:0] hitRefillFlag = _T_303 | _T_310; // @[EmbeddedTLB.scala 222:69]
  wire [39:0] _T_313 = {10'h0,hitData_ppn,2'h0,hitRefillFlag}; // @[Cat.scala 29:58]
  reg [39:0] hitWBStore; // @[Reg.scala 15:16]
  wire  hitExec = hitCheck & hitFlag_x; // @[EmbeddedTLB.scala 227:26]
  reg  _T_327; // @[EmbeddedTLB.scala 236:26]
  reg  _T_328; // @[EmbeddedTLB.scala 237:27]
  reg [63:0] memRespStore; // @[EmbeddedTLB.scala 250:25]
  reg [17:0] missMaskStore; // @[EmbeddedTLB.scala 252:26]
  wire [1:0] memRdata_rsw = io_mem_resp_bits_rdata[9:8]; // @[EmbeddedTLB.scala 255:49]
  wire [19:0] memRdata_ppn = io_mem_resp_bits_rdata[29:10]; // @[EmbeddedTLB.scala 255:49]
  wire [33:0] memRdata_reserved = io_mem_resp_bits_rdata[63:30]; // @[EmbeddedTLB.scala 255:49]
  reg [31:0] raddr; // @[EmbeddedTLB.scala 256:18]
  wire  _T_365 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  reg  alreadyOutFire; // @[Reg.scala 27:20]
  wire  _GEN_2 = _T_365 | alreadyOutFire; // @[Reg.scala 28:19]
  wire [31:0] _T_376 = {satp_ppn,vpn_vpn2,3'h0}; // @[Cat.scala 29:58]
  wire  _T_378 = io_mem_req_ready & io_mem_req_valid; // @[Decoupled.scala 40:37]
  reg [63:0] _T_417; // @[GTimer.scala 24:20]
  wire [63:0] _T_419 = _T_417 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_423 = ~reset; // @[Debug.scala 56:24]
  wire [8:0] _T_448 = _T_400 ? vpn_vpn1 : vpn_vpn0; // @[EmbeddedTLB.scala 311:50]
  wire [31:0] _T_450 = {memRdata_ppn,_T_448,3'h0}; // @[Cat.scala 29:58]
  wire [63:0] _T_472 = {56'h0,io_in_bits_cmd[0],7'h40}; // @[Cat.scala 29:58]
  wire [7:0] _T_482 = {_T_387[7],_T_387[6],_T_387[5],_T_387[4],_T_387[3],_T_387[2],_T_387[1],_T_387[0]}; // @[EmbeddedTLB.scala 320:79]
  wire [7:0] _T_483 = _T_303 | _T_482; // @[EmbeddedTLB.scala 320:68]
  wire [63:0] _T_484 = io_mem_resp_bits_rdata | _T_472; // @[EmbeddedTLB.scala 321:50]
  wire  _GEN_25 = _T_495 ? 1'h0 : 1'h1; // @[EmbeddedTLB.scala 330:80]
  wire [17:0] _T_508 = _T_401 ? 18'h3fe00 : 18'h3ffff; // @[EmbeddedTLB.scala 339:59]
  wire [17:0] _T_509 = _T_400 ? 18'h0 : _T_508; // @[EmbeddedTLB.scala 339:26]
  wire [7:0] _GEN_26 = _T_451 ? _T_483 : 8'h0; // @[EmbeddedTLB.scala 313:36]
  wire  _GEN_31 = _T_451 & _GEN_25; // @[EmbeddedTLB.scala 313:36]
  wire [17:0] _GEN_32 = _T_451 ? _T_509 : 18'h3ffff; // @[EmbeddedTLB.scala 313:36]
  wire [17:0] _GEN_41 = _T_403 ? 18'h3ffff : _GEN_32; // @[EmbeddedTLB.scala 297:82]
  wire [17:0] _GEN_60 = _T_397 ? _GEN_41 : 18'h3ffff; // @[EmbeddedTLB.scala 293:33]
  wire [17:0] _GEN_84 = _T_379 ? _GEN_60 : 18'h3ffff; // @[Conditional.scala 39:67]
  wire [17:0] _GEN_97 = _T_377 ? 18'h3ffff : _GEN_84; // @[Conditional.scala 39:67]
  wire [17:0] missMask = _T_370 ? 18'h3ffff : _GEN_97; // @[Conditional.scala 40:58]
  wire [7:0] _GEN_38 = _T_403 ? 8'h0 : _GEN_26; // @[EmbeddedTLB.scala 297:82]
  wire  _GEN_40 = _T_403 ? 1'h0 : _GEN_31; // @[EmbeddedTLB.scala 297:82]
  wire [1:0] _T_511 = level - 2'h1; // @[EmbeddedTLB.scala 342:24]
  wire [7:0] _GEN_57 = _T_397 ? _GEN_38 : 8'h0; // @[EmbeddedTLB.scala 293:33]
  wire  _GEN_59 = _T_397 & _GEN_40; // @[EmbeddedTLB.scala 293:33]
  wire  _T_512 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_514 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_518 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire [7:0] _GEN_81 = _T_379 ? _GEN_57 : 8'h0; // @[Conditional.scala 39:67]
  wire  _GEN_83 = _T_379 & _GEN_59; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_94 = _T_377 ? 8'h0 : _GEN_81; // @[Conditional.scala 39:67]
  wire  _GEN_96 = _T_377 ? 1'h0 : _GEN_83; // @[Conditional.scala 39:67]
  wire [7:0] missRefillFlag = _T_370 ? 8'h0 : _GEN_94; // @[Conditional.scala 40:58]
  wire  missMetaRefill = _T_370 ? 1'h0 : _GEN_96; // @[Conditional.scala 40:58]
  wire  cmd = state == 3'h3; // @[EmbeddedTLB.scala 365:23]
  wire  _T_522 = state == 3'h1; // @[EmbeddedTLB.scala 367:31]
  wire  _T_529 = state == 3'h0; // @[EmbeddedTLB.scala 371:82]
  wire  _T_530 = hitWB & _T_529; // @[EmbeddedTLB.scala 371:73]
  wire  _T_533 = missMetaRefill | _T_530; // @[EmbeddedTLB.scala 371:63]
  reg  _T_534; // @[EmbeddedTLB.scala 371:33]
  reg [3:0] _T_540; // @[EmbeddedTLB.scala 372:21]
  reg [3:0] _T_541; // @[EmbeddedTLB.scala 372:60]
  reg [26:0] _T_544; // @[EmbeddedTLB.scala 372:84]
  reg [15:0] _T_546; // @[EmbeddedTLB.scala 373:19]
  reg [17:0] _T_548; // @[EmbeddedTLB.scala 373:72]
  reg [7:0] _T_550; // @[EmbeddedTLB.scala 374:19]
  reg [19:0] _T_552; // @[EmbeddedTLB.scala 374:77]
  reg [31:0] _T_554; // @[EmbeddedTLB.scala 375:22]
  wire [59:0] _T_556 = {_T_550,_T_552,_T_554}; // @[Cat.scala 29:58]
  wire [60:0] _T_558 = {_T_544,_T_546,_T_548}; // @[Cat.scala 29:58]
  wire [31:0] _T_561 = {hitData_ppn,12'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_564 = {2'h3,hitMeta_mask,12'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_565 = _T_561 & _T_564; // @[BitUtils.scala 32:13]
  wire [31:0] _T_566 = ~_T_564; // @[BitUtils.scala 32:38]
  wire [31:0] _T_567 = io_in_bits_addr[31:0] & _T_566; // @[BitUtils.scala 32:36]
  wire [31:0] _T_568 = _T_565 | _T_567; // @[BitUtils.scala 32:25]
  wire [31:0] _T_583 = {memRespStore[29:10],12'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_586 = {2'h3,missMaskStore,12'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_587 = _T_583 & _T_586; // @[BitUtils.scala 32:13]
  wire [31:0] _T_588 = ~_T_586; // @[BitUtils.scala 32:38]
  wire [31:0] _T_589 = io_in_bits_addr[31:0] & _T_588; // @[BitUtils.scala 32:36]
  wire [31:0] _T_590 = _T_587 | _T_589; // @[BitUtils.scala 32:25]
  wire  _T_592 = ~hitWB; // @[EmbeddedTLB.scala 380:45]
  wire  _T_593 = hit & _T_592; // @[EmbeddedTLB.scala 380:42]
  wire  _T_595 = _T_298 | loadPF; // @[EmbeddedTLB.scala 380:68]
  wire  _T_596 = _T_595 | storePF; // @[EmbeddedTLB.scala 380:78]
  wire  _T_597 = ~_T_596; // @[EmbeddedTLB.scala 380:53]
  wire  _T_598 = state == 3'h4; // @[EmbeddedTLB.scala 380:97]
  wire  _T_599 = _T_593 ? _T_597 : _T_598; // @[EmbeddedTLB.scala 380:37]
  wire  _T_602 = io_out_ready & _T_529; // @[EmbeddedTLB.scala 382:31]
  wire  _T_603 = ~miss; // @[EmbeddedTLB.scala 382:56]
  wire  _T_604 = _T_602 & _T_603; // @[EmbeddedTLB.scala 382:53]
  wire  _T_606 = _T_604 & _T_592; // @[EmbeddedTLB.scala 382:62]
  wire  _T_607 = _T_606 & io_mdReady; // @[EmbeddedTLB.scala 382:72]
  wire  _T_609 = ~_T_298; // @[EmbeddedTLB.scala 382:90]
  wire  _T_610 = ~loadPF; // @[EmbeddedTLB.scala 382:107]
  wire  _T_611 = _T_609 & _T_610; // @[EmbeddedTLB.scala 382:104]
  wire  _T_612 = ~storePF; // @[EmbeddedTLB.scala 382:118]
  wire  _T_613 = _T_611 & _T_612; // @[EmbeddedTLB.scala 382:115]
  reg [63:0] _T_619; // @[GTimer.scala 24:20]
  wire [63:0] _T_621 = _T_619 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_628; // @[GTimer.scala 24:20]
  wire [63:0] _T_630 = _T_628 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_644; // @[GTimer.scala 24:20]
  wire [63:0] _T_646 = _T_644 + 64'h1; // @[GTimer.scala 25:12]
  wire [4:0] _T_656 = {memRdata_flag_u,memRdata_flag_x,memRdata_flag_w,memRdata_flag_r,memRdata_flag_v}; // @[EmbeddedTLB.scala 390:145]
  wire [63:0] _T_662 = {memRdata_reserved,memRdata_ppn,memRdata_rsw,memRdata_flag_d,memRdata_flag_a,memRdata_flag_g,_T_656}; // @[EmbeddedTLB.scala 390:145]
  reg [63:0] _T_663; // @[GTimer.scala 24:20]
  wire [63:0] _T_665 = _T_663 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_768; // @[GTimer.scala 24:20]
  wire [63:0] _T_770 = _T_768 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_833; // @[GTimer.scala 24:20]
  wire [63:0] _T_835 = _T_833 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_842; // @[GTimer.scala 24:20]
  wire [63:0] _T_844 = _T_842 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_851; // @[GTimer.scala 24:20]
  wire [63:0] _T_853 = _T_851 + 64'h1; // @[GTimer.scala 25:12]
  wire  _GEN_116 = ~_T_370; // @[Debug.scala 56:24]
  wire  _GEN_117 = ~_T_377; // @[Debug.scala 56:24]
  wire  _GEN_118 = _GEN_116 & _GEN_117; // @[Debug.scala 56:24]
  wire  _GEN_119 = _GEN_118 & _T_379; // @[Debug.scala 56:24]
  wire  _GEN_120 = _GEN_119 & _T_397; // @[Debug.scala 56:24]
  wire  _GEN_121 = _GEN_120 & _T_403; // @[Debug.scala 56:24]
  wire  _GEN_122 = _GEN_121 & _T_407; // @[Debug.scala 56:24]
  wire  _GEN_123 = _GEN_122 & DISPLAY_ENABLE; // @[Debug.scala 56:24]
  assign io_in_ready = _T_607 & _T_613; // @[EmbeddedTLB.scala 382:15]
  assign io_out_valid = io_in_valid & _T_599; // @[EmbeddedTLB.scala 380:16]
  assign io_out_bits_addr = hit ? _T_568 : _T_590; // @[EmbeddedTLB.scala 378:15 EmbeddedTLB.scala 379:20]
  assign io_out_bits_size = io_in_bits_size; // @[EmbeddedTLB.scala 378:15]
  assign io_out_bits_cmd = io_in_bits_cmd; // @[EmbeddedTLB.scala 378:15]
  assign io_out_bits_wmask = io_in_bits_wmask; // @[EmbeddedTLB.scala 378:15]
  assign io_out_bits_wdata = io_in_bits_wdata; // @[EmbeddedTLB.scala 378:15]
  assign io_mdWrite_wen = _T_534; // @[TLB.scala 214:14]
  assign io_mdWrite_windex = _T_540; // @[TLB.scala 215:17]
  assign io_mdWrite_waymask = _T_541; // @[TLB.scala 216:18]
  assign io_mdWrite_wdata = {_T_558,_T_556}; // @[TLB.scala 217:16]
  assign io_mem_req_valid = _T_522 | cmd; // @[EmbeddedTLB.scala 367:20]
  assign io_mem_req_bits_addr = hitWB ? hitData_pteaddr : raddr; // @[SimpleBus.scala 64:15]
  assign io_mem_req_bits_size = 3'h3; // @[SimpleBus.scala 66:15]
  assign io_mem_req_bits_cmd = {{3'd0}, cmd}; // @[SimpleBus.scala 65:14]
  assign io_mem_req_bits_wmask = 8'hff; // @[SimpleBus.scala 68:16]
  assign io_mem_req_bits_wdata = hitWB ? {{24'd0}, hitWBStore} : memRespStore; // @[SimpleBus.scala 67:16]
  assign io_mem_resp_ready = 1'h1; // @[EmbeddedTLB.scala 368:21]
  assign io_pf_loadPF = _T_327; // @[EmbeddedTLB.scala 199:13 EmbeddedTLB.scala 236:16]
  assign io_pf_storePF = _T_328; // @[EmbeddedTLB.scala 200:14 EmbeddedTLB.scala 237:17]
  assign io_pf_addr = io_in_bits_addr; // @[EmbeddedTLB.scala 201:11]
  assign io_ipf = 1'h0; // @[EmbeddedTLB.scala 384:10]
  assign io_isFinish = _T_365 | _T_298; // @[EmbeddedTLB.scala 385:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  _T_227 = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  level = _RAND_2[1:0];
  _RAND_3 = {2{`RANDOM}};
  hitWBStore = _RAND_3[39:0];
  _RAND_4 = {1{`RANDOM}};
  _T_327 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _T_328 = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  memRespStore = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  missMaskStore = _RAND_7[17:0];
  _RAND_8 = {1{`RANDOM}};
  raddr = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  alreadyOutFire = _RAND_9[0:0];
  _RAND_10 = {2{`RANDOM}};
  _T_417 = _RAND_10[63:0];
  _RAND_11 = {1{`RANDOM}};
  _T_534 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _T_540 = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  _T_541 = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  _T_544 = _RAND_14[26:0];
  _RAND_15 = {1{`RANDOM}};
  _T_546 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  _T_548 = _RAND_16[17:0];
  _RAND_17 = {1{`RANDOM}};
  _T_550 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  _T_552 = _RAND_18[19:0];
  _RAND_19 = {1{`RANDOM}};
  _T_554 = _RAND_19[31:0];
  _RAND_20 = {2{`RANDOM}};
  _T_619 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  _T_628 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  _T_644 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  _T_663 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  _T_768 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  _T_833 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  _T_842 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  _T_851 = _RAND_27[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_227 <= 64'h1234567887654321;
    end else if (_T_235) begin
      _T_227 <= 64'h1;
    end else begin
      _T_227 <= _T_237;
    end
    if (reset) begin
      state <= 3'h0;
    end else if (_T_370) begin
      if (hitWB) begin
        state <= 3'h3;
      end else if (miss) begin
        state <= 3'h1;
      end
    end else if (_T_377) begin
      if (_T_378) begin
        state <= 3'h2;
      end
    end else if (_T_379) begin
      if (_T_397) begin
        if (_T_403) begin
          if (_T_407) begin
            state <= 3'h5;
          end else begin
            state <= 3'h1;
          end
        end else if (_T_451) begin
          if (_T_495) begin
            state <= 3'h5;
          end else begin
            state <= 3'h4;
          end
        end
      end
    end else if (_T_512) begin
      if (_T_378) begin
        state <= 3'h4;
      end
    end else if (_T_514) begin
      if (_GEN_2) begin
        state <= 3'h0;
      end
    end else if (_T_518) begin
      state <= 3'h0;
    end
    if (reset) begin
      level <= 2'h3;
    end else if (_T_370) begin
      if (!(hitWB)) begin
        if (miss) begin
          level <= 2'h3;
        end
      end
    end else if (!(_T_377)) begin
      if (_T_379) begin
        if (_T_397) begin
          level <= _T_511;
        end
      end
    end
    if (hitWB) begin
      hitWBStore <= _T_313;
    end
    if (reset) begin
      _T_327 <= 1'h0;
    end else if (_T_370) begin
      _T_327 <= _T_338;
    end else if (_T_377) begin
      _T_327 <= _T_338;
    end else if (_T_379) begin
      if (_T_397) begin
        if (_T_403) begin
          if (_T_407) begin
            _T_327 <= _T_414;
          end else begin
            _T_327 <= _T_338;
          end
        end else if (_T_451) begin
          if (_T_495) begin
            _T_327 <= _T_414;
          end else begin
            _T_327 <= _T_338;
          end
        end else begin
          _T_327 <= _T_338;
        end
      end else begin
        _T_327 <= _T_338;
      end
    end else begin
      _T_327 <= _T_338;
    end
    if (reset) begin
      _T_328 <= 1'h0;
    end else if (_T_370) begin
      _T_328 <= _T_352;
    end else if (_T_377) begin
      _T_328 <= _T_352;
    end else if (_T_379) begin
      if (_T_397) begin
        if (_T_403) begin
          if (_T_407) begin
            _T_328 <= _T_416;
          end else begin
            _T_328 <= _T_352;
          end
        end else if (_T_451) begin
          if (_T_495) begin
            _T_328 <= _T_416;
          end else begin
            _T_328 <= _T_352;
          end
        end else begin
          _T_328 <= _T_352;
        end
      end else begin
        _T_328 <= _T_352;
      end
    end else begin
      _T_328 <= _T_352;
    end
    if (!(_T_370)) begin
      if (!(_T_377)) begin
        if (_T_379) begin
          if (_T_397) begin
            if (!(_T_403)) begin
              if (_T_451) begin
                memRespStore <= _T_484;
              end
            end
          end
        end
      end
    end
    if (!(_T_370)) begin
      if (!(_T_377)) begin
        if (_T_379) begin
          if (_T_397) begin
            if (!(_T_403)) begin
              if (_T_451) begin
                if (_T_370) begin
                  missMaskStore <= 18'h3ffff;
                end else if (_T_377) begin
                  missMaskStore <= 18'h3ffff;
                end else if (_T_379) begin
                  if (_T_397) begin
                    if (_T_403) begin
                      missMaskStore <= 18'h3ffff;
                    end else if (_T_451) begin
                      if (_T_400) begin
                        missMaskStore <= 18'h0;
                      end else if (_T_401) begin
                        missMaskStore <= 18'h3fe00;
                      end else begin
                        missMaskStore <= 18'h3ffff;
                      end
                    end else begin
                      missMaskStore <= 18'h3ffff;
                    end
                  end else begin
                    missMaskStore <= 18'h3ffff;
                  end
                end else begin
                  missMaskStore <= 18'h3ffff;
                end
              end
            end
          end
        end
      end
    end
    if (_T_370) begin
      if (!(hitWB)) begin
        if (miss) begin
          raddr <= _T_376;
        end
      end
    end else if (!(_T_377)) begin
      if (_T_379) begin
        if (_T_397) begin
          if (_T_403) begin
            if (!(_T_407)) begin
              raddr <= _T_450;
            end
          end
        end
      end
    end
    if (reset) begin
      alreadyOutFire <= 1'h0;
    end else if (_T_370) begin
      if (hitWB) begin
        alreadyOutFire <= 1'h0;
      end else if (miss) begin
        alreadyOutFire <= 1'h0;
      end else begin
        alreadyOutFire <= _GEN_2;
      end
    end else if (_T_377) begin
      alreadyOutFire <= _GEN_2;
    end else if (_T_379) begin
      alreadyOutFire <= _GEN_2;
    end else if (_T_512) begin
      alreadyOutFire <= _GEN_2;
    end else if (_T_514) begin
      if (_GEN_2) begin
        alreadyOutFire <= 1'h0;
      end else begin
        alreadyOutFire <= _GEN_2;
      end
    end else begin
      alreadyOutFire <= _GEN_2;
    end
    if (reset) begin
      _T_417 <= 64'h0;
    end else begin
      _T_417 <= _T_419;
    end
    if (reset) begin
      _T_534 <= 1'h0;
    end else begin
      _T_534 <= _T_533;
    end
    _T_540 <= io_in_bits_addr[15:12];
    if (hit) begin
      _T_541 <= hitVec;
    end else begin
      _T_541 <= victimWaymask;
    end
    _T_544 <= {_T_57,vpn_vpn0};
    if (hitWB) begin
      _T_546 <= hitMeta_asid;
    end else begin
      _T_546 <= satp_asid;
    end
    if (hitWB) begin
      _T_548 <= hitMeta_mask;
    end else if (_T_370) begin
      _T_548 <= 18'h3ffff;
    end else if (_T_377) begin
      _T_548 <= 18'h3ffff;
    end else if (_T_379) begin
      if (_T_397) begin
        if (_T_403) begin
          _T_548 <= 18'h3ffff;
        end else if (_T_451) begin
          if (_T_400) begin
            _T_548 <= 18'h0;
          end else if (_T_401) begin
            _T_548 <= 18'h3fe00;
          end else begin
            _T_548 <= 18'h3ffff;
          end
        end else begin
          _T_548 <= 18'h3ffff;
        end
      end else begin
        _T_548 <= 18'h3ffff;
      end
    end else begin
      _T_548 <= 18'h3ffff;
    end
    if (hitWB) begin
      _T_550 <= hitRefillFlag;
    end else if (_T_370) begin
      _T_550 <= 8'h0;
    end else if (_T_377) begin
      _T_550 <= 8'h0;
    end else if (_T_379) begin
      if (_T_397) begin
        if (_T_403) begin
          _T_550 <= 8'h0;
        end else if (_T_451) begin
          _T_550 <= _T_483;
        end else begin
          _T_550 <= 8'h0;
        end
      end else begin
        _T_550 <= 8'h0;
      end
    end else begin
      _T_550 <= 8'h0;
    end
    if (hitWB) begin
      _T_552 <= hitData_ppn;
    end else begin
      _T_552 <= memRdata_ppn;
    end
    if (hitWB) begin
      _T_554 <= hitData_pteaddr;
    end else begin
      _T_554 <= raddr;
    end
    if (reset) begin
      _T_619 <= 64'h0;
    end else begin
      _T_619 <= _T_621;
    end
    if (reset) begin
      _T_628 <= 64'h0;
    end else begin
      _T_628 <= _T_630;
    end
    if (reset) begin
      _T_644 <= 64'h0;
    end else begin
      _T_644 <= _T_646;
    end
    if (reset) begin
      _T_663 <= 64'h0;
    end else begin
      _T_663 <= _T_665;
    end
    if (reset) begin
      _T_768 <= 64'h0;
    end else begin
      _T_768 <= _T_770;
    end
    if (reset) begin
      _T_833 <= 64'h0;
    end else begin
      _T_833 <= _T_835;
    end
    if (reset) begin
      _T_842 <= 64'h0;
    end else begin
      _T_842 <= _T_844;
    end
    if (reset) begin
      _T_851 <= 64'h0;
    end else begin
      _T_851 <= _T_853;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_423) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec_1: ",_T_417); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_423) begin
          $fwrite(32'h80000002,"tlbException!!! "); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_423) begin
          $fwrite(32'h80000002," req:addr = 0x%x, cmd = %d, size = %d, wmask = 0x%x, wdata = 0x%x  Memreq:DecoupledIO(ready -> %d, valid -> %d, bits -> addr = 0x%x, cmd = %d, size = %d, wmask = 0x%x, wdata = 0x%x)  MemResp:DecoupledIO(ready -> %d, valid -> %d, bits -> rdata = %x, cmd = %d)",io_in_bits_addr,io_in_bits_cmd,io_in_bits_size,io_in_bits_wmask,io_in_bits_wdata,io_mem_req_ready,io_mem_req_valid,io_mem_req_bits_addr,io_mem_req_bits_cmd,io_mem_req_bits_size,io_mem_req_bits_wmask,io_mem_req_bits_wdata,io_mem_resp_ready,io_mem_resp_valid,io_mem_resp_bits_rdata,io_mem_resp_bits_cmd); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_423) begin
          $fwrite(32'h80000002," level:%d",level); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_123 & _T_423) begin
          $fwrite(32'h80000002,"\n"); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_423) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec_1: ",_T_619); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_423) begin
          $fwrite(32'h80000002,"In(%d, %d) Out(%d, %d) InAddr:%x OutAddr:%x cmd:%d \n",io_in_valid,io_in_ready,io_out_valid,io_out_ready,io_in_bits_addr,io_out_bits_addr,io_in_bits_cmd); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_423) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec_1: ",_T_628); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_423) begin
          $fwrite(32'h80000002,"isAMO:%d io.Flush:%d needFlush:%d alreadyOutFire:%d isFinish:%d\n",ISAMO,1'h0,1'h0,alreadyOutFire,io_isFinish); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_423) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec_1: ",_T_644); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_423) begin
          $fwrite(32'h80000002,"hit:%d hitWB:%d hitVPN:%x hitFlag:%x hitPPN:%x hitRefillFlag:%x hitWBStore:%x hitCheck:%d hitExec:%d hitLoad:%d hitStore:%d\n",hit,hitWB,hitMeta_vpn,_T_310,hitData_ppn,hitRefillFlag,hitWBStore,hitCheck,hitExec,hitLoad,hitStore); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_423) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec_1: ",_T_663); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_423) begin
          $fwrite(32'h80000002,"miss:%d state:%d level:%d raddr:%x memRdata:%x missMask:%x missRefillFlag:%x missMetaRefill:%d\n",miss,state,level,raddr,_T_662,missMask,missRefillFlag,missMetaRefill); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_423) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec_1: ",_T_768); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_423) begin
          $fwrite(32'h80000002,"meta/data: (0)%x|%b|%x (1)%x|%b|%x (2)%x|%b|%x (3)%x|%b|%x rread:%d\n",io_md_0[120:94],io_md_0[59:52],io_md_0[51:32],io_md_1[120:94],io_md_1[59:52],io_md_1[51:32],io_md_2[120:94],io_md_2[59:52],io_md_2[51:32],io_md_3[120:94],io_md_3[59:52],io_md_3[51:32],io_mdReady); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_423) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec_1: ",_T_833); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_423) begin
          $fwrite(32'h80000002,"md: wen:%d windex:%x waymask:%x vpn:%x asid:%x mask:%x flag:%x asid:%x ppn:%x pteaddr:%x\n",io_mdWrite_wen,io_mdWrite_windex,io_mdWrite_waymask,io_mdWrite_wdata[120:94],io_mdWrite_wdata[93:78],io_mdWrite_wdata[77:60],io_mdWrite_wdata[59:52],io_mdWrite_wdata[93:78],io_mdWrite_wdata[51:32],io_mdWrite_wdata[31:0]); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_423) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec_1: ",_T_842); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_423) begin
          $fwrite(32'h80000002,"MemReq(%d, %d) MemResp(%d, %d) addr:%x cmd:%d rdata:%x cmd:%d\n",io_mem_req_valid,io_mem_req_ready,io_mem_resp_valid,io_mem_resp_ready,io_mem_req_bits_addr,io_mem_req_bits_cmd,io_mem_resp_bits_rdata,io_mem_resp_bits_cmd); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_423) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLBExec_1: ",_T_851); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_423) begin
          $fwrite(32'h80000002,"io.ipf:%d hitinstrPF:%d missIPF:%d pf.loadPF:%d pf.storePF:%d loadPF:%d storePF:%d\n",io_ipf,1'h0,1'h0,io_pf_loadPF,io_pf_storePF,loadPF,storePF); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module EmbeddedTLBEmpty_1(
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [2:0]  io_in_bits_size,
  input  [3:0]  io_in_bits_cmd,
  input  [7:0]  io_in_bits_wmask,
  input  [63:0] io_in_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [2:0]  io_out_bits_size,
  output [3:0]  io_out_bits_cmd,
  output [7:0]  io_out_bits_wmask,
  output [63:0] io_out_bits_wdata
);
  assign io_in_ready = io_out_ready; // @[EmbeddedTLB.scala 403:10]
  assign io_out_valid = io_in_valid; // @[EmbeddedTLB.scala 403:10]
  assign io_out_bits_addr = io_in_bits_addr; // @[EmbeddedTLB.scala 403:10]
  assign io_out_bits_size = io_in_bits_size; // @[EmbeddedTLB.scala 403:10]
  assign io_out_bits_cmd = io_in_bits_cmd; // @[EmbeddedTLB.scala 403:10]
  assign io_out_bits_wmask = io_in_bits_wmask; // @[EmbeddedTLB.scala 403:10]
  assign io_out_bits_wdata = io_in_bits_wdata; // @[EmbeddedTLB.scala 403:10]
endmodule
module EmbeddedTLBMD_1(
  input          clock,
  input          reset,
  output [120:0] io_tlbmd_0,
  output [120:0] io_tlbmd_1,
  output [120:0] io_tlbmd_2,
  output [120:0] io_tlbmd_3,
  input          io_write_wen,
  input  [3:0]   io_write_windex,
  input  [3:0]   io_write_waymask,
  input  [120:0] io_write_wdata,
  input  [3:0]   io_rindex,
  output         io_ready
);
`ifdef RANDOMIZE_MEM_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [120:0] tlbmd_0 [0:15]; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_0__T_data; // @[EmbeddedTLB.scala 38:18]
  wire [3:0] tlbmd_0__T_addr; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_0__T_9_data; // @[EmbeddedTLB.scala 38:18]
  wire [3:0] tlbmd_0__T_9_addr; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_0__T_9_mask; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_0__T_9_en; // @[EmbeddedTLB.scala 38:18]
  reg [120:0] tlbmd_1 [0:15]; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_1__T_data; // @[EmbeddedTLB.scala 38:18]
  wire [3:0] tlbmd_1__T_addr; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_1__T_9_data; // @[EmbeddedTLB.scala 38:18]
  wire [3:0] tlbmd_1__T_9_addr; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_1__T_9_mask; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_1__T_9_en; // @[EmbeddedTLB.scala 38:18]
  reg [120:0] tlbmd_2 [0:15]; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_2__T_data; // @[EmbeddedTLB.scala 38:18]
  wire [3:0] tlbmd_2__T_addr; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_2__T_9_data; // @[EmbeddedTLB.scala 38:18]
  wire [3:0] tlbmd_2__T_9_addr; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_2__T_9_mask; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_2__T_9_en; // @[EmbeddedTLB.scala 38:18]
  reg [120:0] tlbmd_3 [0:15]; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_3__T_data; // @[EmbeddedTLB.scala 38:18]
  wire [3:0] tlbmd_3__T_addr; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_3__T_9_data; // @[EmbeddedTLB.scala 38:18]
  wire [3:0] tlbmd_3__T_9_addr; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_3__T_9_mask; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_3__T_9_en; // @[EmbeddedTLB.scala 38:18]
  reg  resetState; // @[EmbeddedTLB.scala 42:27]
  reg [3:0] resetSet; // @[Counter.scala 29:33]
  wire  _T_1 = resetSet == 4'hf; // @[Counter.scala 38:24]
  wire [3:0] _T_3 = resetSet + 4'h1; // @[Counter.scala 39:22]
  wire  resetFinish = resetState & _T_1; // @[Counter.scala 67:17]
  wire  _GEN_2 = resetFinish ? 1'h0 : resetState; // @[EmbeddedTLB.scala 44:22]
  wire [3:0] waymask = resetState ? 4'hf : io_write_waymask; // @[EmbeddedTLB.scala 53:20]
  assign tlbmd_0__T_addr = io_rindex;
  assign tlbmd_0__T_data = tlbmd_0[tlbmd_0__T_addr]; // @[EmbeddedTLB.scala 38:18]
  assign tlbmd_0__T_9_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_0__T_9_addr = resetState ? resetSet : io_write_windex;
  assign tlbmd_0__T_9_mask = waymask[0];
  assign tlbmd_0__T_9_en = resetState | io_write_wen;
  assign tlbmd_1__T_addr = io_rindex;
  assign tlbmd_1__T_data = tlbmd_1[tlbmd_1__T_addr]; // @[EmbeddedTLB.scala 38:18]
  assign tlbmd_1__T_9_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_1__T_9_addr = resetState ? resetSet : io_write_windex;
  assign tlbmd_1__T_9_mask = waymask[1];
  assign tlbmd_1__T_9_en = resetState | io_write_wen;
  assign tlbmd_2__T_addr = io_rindex;
  assign tlbmd_2__T_data = tlbmd_2[tlbmd_2__T_addr]; // @[EmbeddedTLB.scala 38:18]
  assign tlbmd_2__T_9_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_2__T_9_addr = resetState ? resetSet : io_write_windex;
  assign tlbmd_2__T_9_mask = waymask[2];
  assign tlbmd_2__T_9_en = resetState | io_write_wen;
  assign tlbmd_3__T_addr = io_rindex;
  assign tlbmd_3__T_data = tlbmd_3[tlbmd_3__T_addr]; // @[EmbeddedTLB.scala 38:18]
  assign tlbmd_3__T_9_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_3__T_9_addr = resetState ? resetSet : io_write_windex;
  assign tlbmd_3__T_9_mask = waymask[3];
  assign tlbmd_3__T_9_en = resetState | io_write_wen;
  assign io_tlbmd_0 = tlbmd_0__T_data; // @[EmbeddedTLB.scala 39:12]
  assign io_tlbmd_1 = tlbmd_1__T_data; // @[EmbeddedTLB.scala 39:12]
  assign io_tlbmd_2 = tlbmd_2__T_data; // @[EmbeddedTLB.scala 39:12]
  assign io_tlbmd_3 = tlbmd_3__T_data; // @[EmbeddedTLB.scala 39:12]
  assign io_ready = ~resetState; // @[EmbeddedTLB.scala 59:12]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {4{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tlbmd_0[initvar] = _RAND_0[120:0];
  _RAND_1 = {4{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tlbmd_1[initvar] = _RAND_1[120:0];
  _RAND_2 = {4{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tlbmd_2[initvar] = _RAND_2[120:0];
  _RAND_3 = {4{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tlbmd_3[initvar] = _RAND_3[120:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  resetState = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  resetSet = _RAND_5[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(tlbmd_0__T_9_en & tlbmd_0__T_9_mask) begin
      tlbmd_0[tlbmd_0__T_9_addr] <= tlbmd_0__T_9_data; // @[EmbeddedTLB.scala 38:18]
    end
    if(tlbmd_1__T_9_en & tlbmd_1__T_9_mask) begin
      tlbmd_1[tlbmd_1__T_9_addr] <= tlbmd_1__T_9_data; // @[EmbeddedTLB.scala 38:18]
    end
    if(tlbmd_2__T_9_en & tlbmd_2__T_9_mask) begin
      tlbmd_2[tlbmd_2__T_9_addr] <= tlbmd_2__T_9_data; // @[EmbeddedTLB.scala 38:18]
    end
    if(tlbmd_3__T_9_en & tlbmd_3__T_9_mask) begin
      tlbmd_3[tlbmd_3__T_9_addr] <= tlbmd_3__T_9_data; // @[EmbeddedTLB.scala 38:18]
    end
    resetState <= reset | _GEN_2;
    if (reset) begin
      resetSet <= 4'h0;
    end else if (resetState) begin
      resetSet <= _T_3;
    end
  end
endmodule
module EmbeddedTLB_1(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [38:0] io_in_req_bits_addr,
  input  [2:0]  io_in_req_bits_size,
  input  [3:0]  io_in_req_bits_cmd,
  input  [7:0]  io_in_req_bits_wmask,
  input  [63:0] io_in_req_bits_wdata,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [2:0]  io_out_req_bits_size,
  output [3:0]  io_out_req_bits_cmd,
  output [7:0]  io_out_req_bits_wmask,
  output [63:0] io_out_req_bits_wdata,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [3:0]  io_out_resp_bits_cmd,
  input  [63:0] io_out_resp_bits_rdata,
  input         io_mem_req_ready,
  output        io_mem_req_valid,
  output [31:0] io_mem_req_bits_addr,
  output [3:0]  io_mem_req_bits_cmd,
  output [63:0] io_mem_req_bits_wdata,
  input         io_mem_resp_valid,
  input  [3:0]  io_mem_resp_bits_cmd,
  input  [63:0] io_mem_resp_bits_rdata,
  input  [1:0]  io_csrMMU_priviledgeMode,
  input         io_csrMMU_status_sum,
  input         io_csrMMU_status_mxr,
  output        io_csrMMU_loadPF,
  output        io_csrMMU_storePF,
  output [38:0] io_csrMMU_addr,
  input         io_cacheEmpty,
  output        io_ipf,
  output        _T_38_0,
  input  [63:0] CSRSATP,
  input         amoReq,
  input         DISPLAY_ENABLE,
  output        vmEnable_0,
  output        _T_37_1,
  input         MOUFlushTLB
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  wire  tlbExec_clock; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_reset; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_in_ready; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_in_valid; // @[EmbeddedTLB.scala 80:23]
  wire [38:0] tlbExec_io_in_bits_addr; // @[EmbeddedTLB.scala 80:23]
  wire [2:0] tlbExec_io_in_bits_size; // @[EmbeddedTLB.scala 80:23]
  wire [3:0] tlbExec_io_in_bits_cmd; // @[EmbeddedTLB.scala 80:23]
  wire [7:0] tlbExec_io_in_bits_wmask; // @[EmbeddedTLB.scala 80:23]
  wire [63:0] tlbExec_io_in_bits_wdata; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_out_ready; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_out_valid; // @[EmbeddedTLB.scala 80:23]
  wire [31:0] tlbExec_io_out_bits_addr; // @[EmbeddedTLB.scala 80:23]
  wire [2:0] tlbExec_io_out_bits_size; // @[EmbeddedTLB.scala 80:23]
  wire [3:0] tlbExec_io_out_bits_cmd; // @[EmbeddedTLB.scala 80:23]
  wire [7:0] tlbExec_io_out_bits_wmask; // @[EmbeddedTLB.scala 80:23]
  wire [63:0] tlbExec_io_out_bits_wdata; // @[EmbeddedTLB.scala 80:23]
  wire [120:0] tlbExec_io_md_0; // @[EmbeddedTLB.scala 80:23]
  wire [120:0] tlbExec_io_md_1; // @[EmbeddedTLB.scala 80:23]
  wire [120:0] tlbExec_io_md_2; // @[EmbeddedTLB.scala 80:23]
  wire [120:0] tlbExec_io_md_3; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mdWrite_wen; // @[EmbeddedTLB.scala 80:23]
  wire [3:0] tlbExec_io_mdWrite_windex; // @[EmbeddedTLB.scala 80:23]
  wire [3:0] tlbExec_io_mdWrite_waymask; // @[EmbeddedTLB.scala 80:23]
  wire [120:0] tlbExec_io_mdWrite_wdata; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mdReady; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mem_req_ready; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mem_req_valid; // @[EmbeddedTLB.scala 80:23]
  wire [31:0] tlbExec_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 80:23]
  wire [2:0] tlbExec_io_mem_req_bits_size; // @[EmbeddedTLB.scala 80:23]
  wire [3:0] tlbExec_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 80:23]
  wire [7:0] tlbExec_io_mem_req_bits_wmask; // @[EmbeddedTLB.scala 80:23]
  wire [63:0] tlbExec_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mem_resp_ready; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mem_resp_valid; // @[EmbeddedTLB.scala 80:23]
  wire [3:0] tlbExec_io_mem_resp_bits_cmd; // @[EmbeddedTLB.scala 80:23]
  wire [63:0] tlbExec_io_mem_resp_bits_rdata; // @[EmbeddedTLB.scala 80:23]
  wire [63:0] tlbExec_io_satp; // @[EmbeddedTLB.scala 80:23]
  wire [1:0] tlbExec_io_pf_priviledgeMode; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_pf_status_sum; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_pf_status_mxr; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_pf_loadPF; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_pf_storePF; // @[EmbeddedTLB.scala 80:23]
  wire [38:0] tlbExec_io_pf_addr; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_ipf; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_isFinish; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_ISAMO; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_DISPLAY_ENABLE; // @[EmbeddedTLB.scala 80:23]
  wire  tlbEmpty_io_in_ready; // @[EmbeddedTLB.scala 81:24]
  wire  tlbEmpty_io_in_valid; // @[EmbeddedTLB.scala 81:24]
  wire [31:0] tlbEmpty_io_in_bits_addr; // @[EmbeddedTLB.scala 81:24]
  wire [2:0] tlbEmpty_io_in_bits_size; // @[EmbeddedTLB.scala 81:24]
  wire [3:0] tlbEmpty_io_in_bits_cmd; // @[EmbeddedTLB.scala 81:24]
  wire [7:0] tlbEmpty_io_in_bits_wmask; // @[EmbeddedTLB.scala 81:24]
  wire [63:0] tlbEmpty_io_in_bits_wdata; // @[EmbeddedTLB.scala 81:24]
  wire  tlbEmpty_io_out_ready; // @[EmbeddedTLB.scala 81:24]
  wire  tlbEmpty_io_out_valid; // @[EmbeddedTLB.scala 81:24]
  wire [31:0] tlbEmpty_io_out_bits_addr; // @[EmbeddedTLB.scala 81:24]
  wire [2:0] tlbEmpty_io_out_bits_size; // @[EmbeddedTLB.scala 81:24]
  wire [3:0] tlbEmpty_io_out_bits_cmd; // @[EmbeddedTLB.scala 81:24]
  wire [7:0] tlbEmpty_io_out_bits_wmask; // @[EmbeddedTLB.scala 81:24]
  wire [63:0] tlbEmpty_io_out_bits_wdata; // @[EmbeddedTLB.scala 81:24]
  wire  mdTLB_clock; // @[EmbeddedTLB.scala 82:21]
  wire  mdTLB_reset; // @[EmbeddedTLB.scala 82:21]
  wire [120:0] mdTLB_io_tlbmd_0; // @[EmbeddedTLB.scala 82:21]
  wire [120:0] mdTLB_io_tlbmd_1; // @[EmbeddedTLB.scala 82:21]
  wire [120:0] mdTLB_io_tlbmd_2; // @[EmbeddedTLB.scala 82:21]
  wire [120:0] mdTLB_io_tlbmd_3; // @[EmbeddedTLB.scala 82:21]
  wire  mdTLB_io_write_wen; // @[EmbeddedTLB.scala 82:21]
  wire [3:0] mdTLB_io_write_windex; // @[EmbeddedTLB.scala 82:21]
  wire [3:0] mdTLB_io_write_waymask; // @[EmbeddedTLB.scala 82:21]
  wire [120:0] mdTLB_io_write_wdata; // @[EmbeddedTLB.scala 82:21]
  wire [3:0] mdTLB_io_rindex; // @[EmbeddedTLB.scala 82:21]
  wire  mdTLB_io_ready; // @[EmbeddedTLB.scala 82:21]
  reg [120:0] _T__0; // @[Reg.scala 15:16]
  reg [120:0] _T__1; // @[Reg.scala 15:16]
  reg [120:0] _T__2; // @[Reg.scala 15:16]
  reg [120:0] _T__3; // @[Reg.scala 15:16]
  wire  mdUpdate = io_in_req_valid & tlbExec_io_in_ready; // @[EmbeddedTLB.scala 114:26]
  wire  _T_14 = CSRSATP[63:60] == 4'h8; // @[EmbeddedTLB.scala 102:49]
  wire  _T_15 = io_csrMMU_priviledgeMode < 2'h3; // @[EmbeddedTLB.scala 102:86]
  wire  vmEnable = _T_14 & _T_15; // @[EmbeddedTLB.scala 102:57]
  reg  _T_16; // @[EmbeddedTLB.scala 105:24]
  wire  _GEN_4 = tlbExec_io_isFinish ? 1'h0 : _T_16; // @[EmbeddedTLB.scala 106:25]
  wire  _T_18 = mdUpdate & vmEnable; // @[EmbeddedTLB.scala 107:37]
  wire  _GEN_5 = _T_18 | _GEN_4; // @[EmbeddedTLB.scala 107:50]
  reg [38:0] _T_20_addr; // @[Reg.scala 15:16]
  reg [2:0] _T_20_size; // @[Reg.scala 15:16]
  reg [3:0] _T_20_cmd; // @[Reg.scala 15:16]
  reg [7:0] _T_20_wmask; // @[Reg.scala 15:16]
  reg [63:0] _T_20_wdata; // @[Reg.scala 15:16]
  wire  _T_22 = tlbEmpty_io_out_ready & tlbEmpty_io_out_valid; // @[Decoupled.scala 40:37]
  reg  _T_23; // @[Pipeline.scala 24:24]
  wire  _GEN_12 = _T_22 ? 1'h0 : _T_23; // @[Pipeline.scala 25:25]
  wire  _T_24 = tlbExec_io_out_valid & tlbEmpty_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_13 = _T_24 | _GEN_12; // @[Pipeline.scala 26:38]
  reg [31:0] _T_26_addr; // @[Reg.scala 15:16]
  reg [2:0] _T_26_size; // @[Reg.scala 15:16]
  reg [3:0] _T_26_cmd; // @[Reg.scala 15:16]
  reg [7:0] _T_26_wmask; // @[Reg.scala 15:16]
  reg [63:0] _T_26_wdata; // @[Reg.scala 15:16]
  wire  _T_27 = ~vmEnable; // @[EmbeddedTLB.scala 123:8]
  wire  _T_29 = ~tlbExec_io_out_ready; // @[EmbeddedTLB.scala 142:84]
  wire  _T_30 = tlbExec_io_out_valid & _T_29; // @[EmbeddedTLB.scala 142:81]
  reg  _T_31; // @[Reg.scala 27:20]
  wire  _GEN_29 = _T_30 | _T_31; // @[Reg.scala 28:19]
  wire  _T_32 = tlbExec_io_out_ready & tlbExec_io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_33 = _T_31 & _T_32; // @[EmbeddedTLB.scala 143:27]
  wire  _T_34 = ~_T_31; // @[EmbeddedTLB.scala 144:46]
  wire  _T_35 = tlbExec_io_out_valid & _T_34; // @[EmbeddedTLB.scala 144:43]
  wire  _T_36 = tlbExec_io_pf_loadPF | tlbExec_io_pf_storePF; // @[Bundle.scala 135:23]
  wire  _T_37 = _T_35 | _T_36; // @[EmbeddedTLB.scala 144:65]
  wire  _T_38 = io_csrMMU_loadPF | io_csrMMU_storePF; // @[Bundle.scala 135:23]
  reg [63:0] _T_39; // @[GTimer.scala 24:20]
  wire [63:0] _T_41 = _T_39 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_45 = ~reset; // @[Debug.scala 56:24]
  reg [63:0] _T_48; // @[GTimer.scala 24:20]
  wire [63:0] _T_50 = _T_48 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_57; // @[GTimer.scala 24:20]
  wire [63:0] _T_59 = _T_57 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_66; // @[GTimer.scala 24:20]
  wire [63:0] _T_68 = _T_66 + 64'h1; // @[GTimer.scala 25:12]
  EmbeddedTLBExec_1 tlbExec ( // @[EmbeddedTLB.scala 80:23]
    .clock(tlbExec_clock),
    .reset(tlbExec_reset),
    .io_in_ready(tlbExec_io_in_ready),
    .io_in_valid(tlbExec_io_in_valid),
    .io_in_bits_addr(tlbExec_io_in_bits_addr),
    .io_in_bits_size(tlbExec_io_in_bits_size),
    .io_in_bits_cmd(tlbExec_io_in_bits_cmd),
    .io_in_bits_wmask(tlbExec_io_in_bits_wmask),
    .io_in_bits_wdata(tlbExec_io_in_bits_wdata),
    .io_out_ready(tlbExec_io_out_ready),
    .io_out_valid(tlbExec_io_out_valid),
    .io_out_bits_addr(tlbExec_io_out_bits_addr),
    .io_out_bits_size(tlbExec_io_out_bits_size),
    .io_out_bits_cmd(tlbExec_io_out_bits_cmd),
    .io_out_bits_wmask(tlbExec_io_out_bits_wmask),
    .io_out_bits_wdata(tlbExec_io_out_bits_wdata),
    .io_md_0(tlbExec_io_md_0),
    .io_md_1(tlbExec_io_md_1),
    .io_md_2(tlbExec_io_md_2),
    .io_md_3(tlbExec_io_md_3),
    .io_mdWrite_wen(tlbExec_io_mdWrite_wen),
    .io_mdWrite_windex(tlbExec_io_mdWrite_windex),
    .io_mdWrite_waymask(tlbExec_io_mdWrite_waymask),
    .io_mdWrite_wdata(tlbExec_io_mdWrite_wdata),
    .io_mdReady(tlbExec_io_mdReady),
    .io_mem_req_ready(tlbExec_io_mem_req_ready),
    .io_mem_req_valid(tlbExec_io_mem_req_valid),
    .io_mem_req_bits_addr(tlbExec_io_mem_req_bits_addr),
    .io_mem_req_bits_size(tlbExec_io_mem_req_bits_size),
    .io_mem_req_bits_cmd(tlbExec_io_mem_req_bits_cmd),
    .io_mem_req_bits_wmask(tlbExec_io_mem_req_bits_wmask),
    .io_mem_req_bits_wdata(tlbExec_io_mem_req_bits_wdata),
    .io_mem_resp_ready(tlbExec_io_mem_resp_ready),
    .io_mem_resp_valid(tlbExec_io_mem_resp_valid),
    .io_mem_resp_bits_cmd(tlbExec_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_rdata(tlbExec_io_mem_resp_bits_rdata),
    .io_satp(tlbExec_io_satp),
    .io_pf_priviledgeMode(tlbExec_io_pf_priviledgeMode),
    .io_pf_status_sum(tlbExec_io_pf_status_sum),
    .io_pf_status_mxr(tlbExec_io_pf_status_mxr),
    .io_pf_loadPF(tlbExec_io_pf_loadPF),
    .io_pf_storePF(tlbExec_io_pf_storePF),
    .io_pf_addr(tlbExec_io_pf_addr),
    .io_ipf(tlbExec_io_ipf),
    .io_isFinish(tlbExec_io_isFinish),
    .ISAMO(tlbExec_ISAMO),
    .DISPLAY_ENABLE(tlbExec_DISPLAY_ENABLE)
  );
  EmbeddedTLBEmpty_1 tlbEmpty ( // @[EmbeddedTLB.scala 81:24]
    .io_in_ready(tlbEmpty_io_in_ready),
    .io_in_valid(tlbEmpty_io_in_valid),
    .io_in_bits_addr(tlbEmpty_io_in_bits_addr),
    .io_in_bits_size(tlbEmpty_io_in_bits_size),
    .io_in_bits_cmd(tlbEmpty_io_in_bits_cmd),
    .io_in_bits_wmask(tlbEmpty_io_in_bits_wmask),
    .io_in_bits_wdata(tlbEmpty_io_in_bits_wdata),
    .io_out_ready(tlbEmpty_io_out_ready),
    .io_out_valid(tlbEmpty_io_out_valid),
    .io_out_bits_addr(tlbEmpty_io_out_bits_addr),
    .io_out_bits_size(tlbEmpty_io_out_bits_size),
    .io_out_bits_cmd(tlbEmpty_io_out_bits_cmd),
    .io_out_bits_wmask(tlbEmpty_io_out_bits_wmask),
    .io_out_bits_wdata(tlbEmpty_io_out_bits_wdata)
  );
  EmbeddedTLBMD_1 mdTLB ( // @[EmbeddedTLB.scala 82:21]
    .clock(mdTLB_clock),
    .reset(mdTLB_reset),
    .io_tlbmd_0(mdTLB_io_tlbmd_0),
    .io_tlbmd_1(mdTLB_io_tlbmd_1),
    .io_tlbmd_2(mdTLB_io_tlbmd_2),
    .io_tlbmd_3(mdTLB_io_tlbmd_3),
    .io_write_wen(mdTLB_io_write_wen),
    .io_write_windex(mdTLB_io_write_windex),
    .io_write_waymask(mdTLB_io_write_waymask),
    .io_write_wdata(mdTLB_io_write_wdata),
    .io_rindex(mdTLB_io_rindex),
    .io_ready(mdTLB_io_ready)
  );
  assign io_in_req_ready = _T_27 ? io_out_req_ready : tlbExec_io_in_ready; // @[EmbeddedTLB.scala 110:16 EmbeddedTLB.scala 127:21]
  assign io_in_resp_valid = io_out_resp_valid; // @[EmbeddedTLB.scala 138:15]
  assign io_in_resp_bits_cmd = io_out_resp_bits_cmd; // @[EmbeddedTLB.scala 138:15]
  assign io_in_resp_bits_rdata = io_out_resp_bits_rdata; // @[EmbeddedTLB.scala 138:15]
  assign io_out_req_valid = _T_27 ? io_in_req_valid : tlbEmpty_io_out_valid; // @[EmbeddedTLB.scala 126:22 EmbeddedTLB.scala 135:41]
  assign io_out_req_bits_addr = _T_27 ? io_in_req_bits_addr[31:0] : tlbEmpty_io_out_bits_addr; // @[EmbeddedTLB.scala 128:26 EmbeddedTLB.scala 135:41]
  assign io_out_req_bits_size = _T_27 ? io_in_req_bits_size : tlbEmpty_io_out_bits_size; // @[EmbeddedTLB.scala 129:26 EmbeddedTLB.scala 135:41]
  assign io_out_req_bits_cmd = _T_27 ? io_in_req_bits_cmd : tlbEmpty_io_out_bits_cmd; // @[EmbeddedTLB.scala 130:25 EmbeddedTLB.scala 135:41]
  assign io_out_req_bits_wmask = _T_27 ? io_in_req_bits_wmask : tlbEmpty_io_out_bits_wmask; // @[EmbeddedTLB.scala 131:27 EmbeddedTLB.scala 135:41]
  assign io_out_req_bits_wdata = _T_27 ? io_in_req_bits_wdata : tlbEmpty_io_out_bits_wdata; // @[EmbeddedTLB.scala 132:27 EmbeddedTLB.scala 135:41]
  assign io_out_resp_ready = 1'h1; // @[EmbeddedTLB.scala 138:15]
  assign io_mem_req_valid = tlbExec_io_mem_req_valid; // @[EmbeddedTLB.scala 87:18]
  assign io_mem_req_bits_addr = tlbExec_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 87:18]
  assign io_mem_req_bits_cmd = tlbExec_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 87:18]
  assign io_mem_req_bits_wdata = tlbExec_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 87:18]
  assign io_csrMMU_loadPF = tlbExec_io_pf_loadPF; // @[EmbeddedTLB.scala 88:17]
  assign io_csrMMU_storePF = tlbExec_io_pf_storePF; // @[EmbeddedTLB.scala 88:17]
  assign io_csrMMU_addr = tlbExec_io_pf_addr; // @[EmbeddedTLB.scala 88:17]
  assign io_ipf = 1'h0; // @[EmbeddedTLB.scala 94:10]
  assign _T_38_0 = _T_38;
  assign vmEnable_0 = vmEnable;
  assign _T_37_1 = _T_37;
  assign tlbExec_clock = clock;
  assign tlbExec_reset = reset;
  assign tlbExec_io_in_valid = _T_16; // @[EmbeddedTLB.scala 112:17]
  assign tlbExec_io_in_bits_addr = _T_20_addr; // @[EmbeddedTLB.scala 111:16]
  assign tlbExec_io_in_bits_size = _T_20_size; // @[EmbeddedTLB.scala 111:16]
  assign tlbExec_io_in_bits_cmd = _T_20_cmd; // @[EmbeddedTLB.scala 111:16]
  assign tlbExec_io_in_bits_wmask = _T_20_wmask; // @[EmbeddedTLB.scala 111:16]
  assign tlbExec_io_in_bits_wdata = _T_20_wdata; // @[EmbeddedTLB.scala 111:16]
  assign tlbExec_io_out_ready = _T_27 | tlbEmpty_io_in_ready; // @[Pipeline.scala 29:16 EmbeddedTLB.scala 124:26]
  assign tlbExec_io_md_0 = _T__0; // @[EmbeddedTLB.scala 89:17]
  assign tlbExec_io_md_1 = _T__1; // @[EmbeddedTLB.scala 89:17]
  assign tlbExec_io_md_2 = _T__2; // @[EmbeddedTLB.scala 89:17]
  assign tlbExec_io_md_3 = _T__3; // @[EmbeddedTLB.scala 89:17]
  assign tlbExec_io_mdReady = mdTLB_io_ready; // @[EmbeddedTLB.scala 90:22]
  assign tlbExec_io_mem_req_ready = io_mem_req_ready; // @[EmbeddedTLB.scala 87:18]
  assign tlbExec_io_mem_resp_valid = io_mem_resp_valid; // @[EmbeddedTLB.scala 87:18]
  assign tlbExec_io_mem_resp_bits_cmd = io_mem_resp_bits_cmd; // @[EmbeddedTLB.scala 87:18]
  assign tlbExec_io_mem_resp_bits_rdata = io_mem_resp_bits_rdata; // @[EmbeddedTLB.scala 87:18]
  assign tlbExec_io_satp = CSRSATP; // @[EmbeddedTLB.scala 86:19]
  assign tlbExec_io_pf_priviledgeMode = io_csrMMU_priviledgeMode; // @[EmbeddedTLB.scala 88:17]
  assign tlbExec_io_pf_status_sum = io_csrMMU_status_sum; // @[EmbeddedTLB.scala 88:17]
  assign tlbExec_io_pf_status_mxr = io_csrMMU_status_mxr; // @[EmbeddedTLB.scala 88:17]
  assign tlbExec_ISAMO = amoReq;
  assign tlbExec_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign tlbEmpty_io_in_valid = _T_23; // @[Pipeline.scala 31:17]
  assign tlbEmpty_io_in_bits_addr = _T_26_addr; // @[Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_size = _T_26_size; // @[Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_cmd = _T_26_cmd; // @[Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_wmask = _T_26_wmask; // @[Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_wdata = _T_26_wdata; // @[Pipeline.scala 30:16]
  assign tlbEmpty_io_out_ready = _T_27 | io_out_req_ready; // @[EmbeddedTLB.scala 125:52 EmbeddedTLB.scala 135:41]
  assign mdTLB_clock = clock;
  assign mdTLB_reset = reset | MOUFlushTLB; // @[EmbeddedTLB.scala 99:15]
  assign mdTLB_io_write_wen = tlbExec_io_mdWrite_wen; // @[EmbeddedTLB.scala 92:18]
  assign mdTLB_io_write_windex = tlbExec_io_mdWrite_windex; // @[EmbeddedTLB.scala 92:18]
  assign mdTLB_io_write_waymask = tlbExec_io_mdWrite_waymask; // @[EmbeddedTLB.scala 92:18]
  assign mdTLB_io_write_wdata = tlbExec_io_mdWrite_wdata; // @[EmbeddedTLB.scala 92:18]
  assign mdTLB_io_rindex = io_in_req_bits_addr[15:12]; // @[EmbeddedTLB.scala 91:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  _T__0 = _RAND_0[120:0];
  _RAND_1 = {4{`RANDOM}};
  _T__1 = _RAND_1[120:0];
  _RAND_2 = {4{`RANDOM}};
  _T__2 = _RAND_2[120:0];
  _RAND_3 = {4{`RANDOM}};
  _T__3 = _RAND_3[120:0];
  _RAND_4 = {1{`RANDOM}};
  _T_16 = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  _T_20_addr = _RAND_5[38:0];
  _RAND_6 = {1{`RANDOM}};
  _T_20_size = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  _T_20_cmd = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  _T_20_wmask = _RAND_8[7:0];
  _RAND_9 = {2{`RANDOM}};
  _T_20_wdata = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  _T_23 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _T_26_addr = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  _T_26_size = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  _T_26_cmd = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  _T_26_wmask = _RAND_14[7:0];
  _RAND_15 = {2{`RANDOM}};
  _T_26_wdata = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  _T_31 = _RAND_16[0:0];
  _RAND_17 = {2{`RANDOM}};
  _T_39 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  _T_48 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  _T_57 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  _T_66 = _RAND_20[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (mdUpdate) begin
      _T__0 <= mdTLB_io_tlbmd_0;
    end
    if (mdUpdate) begin
      _T__1 <= mdTLB_io_tlbmd_1;
    end
    if (mdUpdate) begin
      _T__2 <= mdTLB_io_tlbmd_2;
    end
    if (mdUpdate) begin
      _T__3 <= mdTLB_io_tlbmd_3;
    end
    if (reset) begin
      _T_16 <= 1'h0;
    end else begin
      _T_16 <= _GEN_5;
    end
    if (mdUpdate) begin
      _T_20_addr <= io_in_req_bits_addr;
    end
    if (mdUpdate) begin
      _T_20_size <= io_in_req_bits_size;
    end
    if (mdUpdate) begin
      _T_20_cmd <= io_in_req_bits_cmd;
    end
    if (mdUpdate) begin
      _T_20_wmask <= io_in_req_bits_wmask;
    end
    if (mdUpdate) begin
      _T_20_wdata <= io_in_req_bits_wdata;
    end
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _GEN_13;
    end
    if (_T_24) begin
      _T_26_addr <= tlbExec_io_out_bits_addr;
    end
    if (_T_24) begin
      _T_26_size <= tlbExec_io_out_bits_size;
    end
    if (_T_24) begin
      _T_26_cmd <= tlbExec_io_out_bits_cmd;
    end
    if (_T_24) begin
      _T_26_wmask <= tlbExec_io_out_bits_wmask;
    end
    if (_T_24) begin
      _T_26_wdata <= tlbExec_io_out_bits_wdata;
    end
    if (reset) begin
      _T_31 <= 1'h0;
    end else if (_T_33) begin
      _T_31 <= 1'h0;
    end else begin
      _T_31 <= _GEN_29;
    end
    if (reset) begin
      _T_39 <= 64'h0;
    end else begin
      _T_39 <= _T_41;
    end
    if (reset) begin
      _T_48 <= 64'h0;
    end else begin
      _T_48 <= _T_50;
    end
    if (reset) begin
      _T_57 <= 64'h0;
    end else begin
      _T_57 <= _T_59;
    end
    if (reset) begin
      _T_66 <= 64'h0;
    end else begin
      _T_66 <= _T_68;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_45) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLB_1: ",_T_39); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_45) begin
          $fwrite(32'h80000002,"InReq(%d, %d) InResp(%d, %d) OutReq(%d, %d) OutResp(%d, %d) vmEnable:%d mode:%d\n",io_in_req_valid,io_in_req_ready,io_in_resp_valid,1'h1,io_out_req_valid,io_out_req_ready,io_out_resp_valid,io_out_resp_ready,vmEnable,io_csrMMU_priviledgeMode); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_45) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLB_1: ",_T_48); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_45) begin
          $fwrite(32'h80000002,"InReq: addr:%x cmd:%d wdata:%x OutReq: addr:%x cmd:%x wdata:%x\n",io_in_req_bits_addr,io_in_req_bits_cmd,io_in_req_bits_wdata,io_out_req_bits_addr,io_out_req_bits_cmd,io_out_req_bits_wdata); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_45) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLB_1: ",_T_57); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_45) begin
          $fwrite(32'h80000002,"OutResp: rdata:%x cmd:%x Inresp: rdata:%x cmd:%x\n",io_out_resp_bits_rdata,io_out_resp_bits_cmd,io_in_resp_bits_rdata,io_in_resp_bits_cmd); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_45) begin
          $fwrite(32'h80000002,"[%d] EmbeddedTLB_1: ",_T_66); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_45) begin
          $fwrite(32'h80000002,"satp:%x flush:%d cacheEmpty:%d instrPF:%d loadPF:%d storePF:%d \n",CSRSATP,1'h0,io_cacheEmpty,io_ipf,io_csrMMU_loadPF,io_csrMMU_storePF); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CacheStage1_1(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [2:0]  io_in_bits_size,
  input  [3:0]  io_in_bits_cmd,
  input  [7:0]  io_in_bits_wmask,
  input  [63:0] io_in_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_req_addr,
  output [2:0]  io_out_bits_req_size,
  output [3:0]  io_out_bits_req_cmd,
  output [7:0]  io_out_bits_req_wmask,
  output [63:0] io_out_bits_req_wdata,
  input         io_metaReadBus_req_ready,
  output        io_metaReadBus_req_valid,
  output [6:0]  io_metaReadBus_req_bits_setIdx,
  input  [18:0] io_metaReadBus_resp_data_0_tag,
  input         io_metaReadBus_resp_data_0_valid,
  input         io_metaReadBus_resp_data_0_dirty,
  input  [18:0] io_metaReadBus_resp_data_1_tag,
  input         io_metaReadBus_resp_data_1_valid,
  input         io_metaReadBus_resp_data_1_dirty,
  input  [18:0] io_metaReadBus_resp_data_2_tag,
  input         io_metaReadBus_resp_data_2_valid,
  input         io_metaReadBus_resp_data_2_dirty,
  input  [18:0] io_metaReadBus_resp_data_3_tag,
  input         io_metaReadBus_resp_data_3_valid,
  input         io_metaReadBus_resp_data_3_dirty,
  input         io_dataReadBus_req_ready,
  output        io_dataReadBus_req_valid,
  output [9:0]  io_dataReadBus_req_bits_setIdx,
  input  [63:0] io_dataReadBus_resp_data_0_data,
  input  [63:0] io_dataReadBus_resp_data_1_data,
  input  [63:0] io_dataReadBus_resp_data_2_data,
  input  [63:0] io_dataReadBus_resp_data_3_data,
  input         DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  _T = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  reg [63:0] _T_1; // @[GTimer.scala 24:20]
  wire [63:0] _T_3 = _T_1 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_5 = _T & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  wire  _T_7 = ~reset; // @[Debug.scala 56:24]
  wire  _T_29 = io_in_valid & io_metaReadBus_req_ready; // @[Cache.scala 133:31]
  wire  _T_31 = ~io_in_valid; // @[Cache.scala 134:19]
  wire  _T_32 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_33 = _T_31 | _T_32; // @[Cache.scala 134:32]
  wire  _T_34 = _T_33 & io_metaReadBus_req_ready; // @[Cache.scala 134:50]
  reg [63:0] _T_36; // @[GTimer.scala 24:20]
  wire [63:0] _T_38 = _T_36 + 64'h1; // @[GTimer.scala 25:12]
  assign io_in_ready = _T_34 & io_dataReadBus_req_ready; // @[Cache.scala 134:15]
  assign io_out_valid = _T_29 & io_dataReadBus_req_ready; // @[Cache.scala 133:16]
  assign io_out_bits_req_addr = io_in_bits_addr; // @[Cache.scala 132:19]
  assign io_out_bits_req_size = io_in_bits_size; // @[Cache.scala 132:19]
  assign io_out_bits_req_cmd = io_in_bits_cmd; // @[Cache.scala 132:19]
  assign io_out_bits_req_wmask = io_in_bits_wmask; // @[Cache.scala 132:19]
  assign io_out_bits_req_wdata = io_in_bits_wdata; // @[Cache.scala 132:19]
  assign io_metaReadBus_req_valid = io_in_valid & io_out_ready; // @[SRAMTemplate.scala 53:20]
  assign io_metaReadBus_req_bits_setIdx = io_in_bits_addr[12:6]; // @[SRAMTemplate.scala 26:17]
  assign io_dataReadBus_req_valid = io_in_valid & io_out_ready; // @[SRAMTemplate.scala 53:20]
  assign io_dataReadBus_req_bits_setIdx = {io_in_bits_addr[12:6],io_in_bits_addr[5:3]}; // @[SRAMTemplate.scala 26:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  _T_1 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  _T_36 = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_1 <= 64'h0;
    end else begin
      _T_1 <= _T_3;
    end
    if (reset) begin
      _T_36 <= 64'h0;
    end else begin
      _T_36 <= _T_38;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5 & _T_7) begin
          $fwrite(32'h80000002,"[%d] CacheStage1_1: ",_T_1); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5 & _T_7) begin
          $fwrite(32'h80000002,"[L1$] cache stage1, addr in: %x, user: %x id: %x\n",io_in_bits_addr,1'h0,1'h0); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_7) begin
          $fwrite(32'h80000002,"[%d] CacheStage1_1: ",_T_36); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_7) begin
          $fwrite(32'h80000002,"in.ready = %d, in.valid = %d, out.valid = %d, out.ready = %d, addr = %x, cmd = %x, dataReadBus.req.valid = %d\n",io_in_ready,io_in_valid,io_out_valid,io_out_ready,io_in_bits_addr,io_in_bits_cmd,io_dataReadBus_req_valid); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CacheStage2_1(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_req_addr,
  input  [2:0]  io_in_bits_req_size,
  input  [3:0]  io_in_bits_req_cmd,
  input  [7:0]  io_in_bits_req_wmask,
  input  [63:0] io_in_bits_req_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_req_addr,
  output [2:0]  io_out_bits_req_size,
  output [3:0]  io_out_bits_req_cmd,
  output [7:0]  io_out_bits_req_wmask,
  output [63:0] io_out_bits_req_wdata,
  output [18:0] io_out_bits_metas_0_tag,
  output        io_out_bits_metas_0_valid,
  output        io_out_bits_metas_0_dirty,
  output [18:0] io_out_bits_metas_1_tag,
  output        io_out_bits_metas_1_valid,
  output        io_out_bits_metas_1_dirty,
  output [18:0] io_out_bits_metas_2_tag,
  output        io_out_bits_metas_2_valid,
  output        io_out_bits_metas_2_dirty,
  output [18:0] io_out_bits_metas_3_tag,
  output        io_out_bits_metas_3_valid,
  output        io_out_bits_metas_3_dirty,
  output [63:0] io_out_bits_datas_0_data,
  output [63:0] io_out_bits_datas_1_data,
  output [63:0] io_out_bits_datas_2_data,
  output [63:0] io_out_bits_datas_3_data,
  output        io_out_bits_hit,
  output [3:0]  io_out_bits_waymask,
  output        io_out_bits_mmio,
  output        io_out_bits_isForwardData,
  output [63:0] io_out_bits_forwardData_data_data,
  output [3:0]  io_out_bits_forwardData_waymask,
  input  [18:0] io_metaReadResp_0_tag,
  input         io_metaReadResp_0_valid,
  input         io_metaReadResp_0_dirty,
  input  [18:0] io_metaReadResp_1_tag,
  input         io_metaReadResp_1_valid,
  input         io_metaReadResp_1_dirty,
  input  [18:0] io_metaReadResp_2_tag,
  input         io_metaReadResp_2_valid,
  input         io_metaReadResp_2_dirty,
  input  [18:0] io_metaReadResp_3_tag,
  input         io_metaReadResp_3_valid,
  input         io_metaReadResp_3_dirty,
  input  [63:0] io_dataReadResp_0_data,
  input  [63:0] io_dataReadResp_1_data,
  input  [63:0] io_dataReadResp_2_data,
  input  [63:0] io_dataReadResp_3_data,
  input         io_metaWriteBus_req_valid,
  input  [6:0]  io_metaWriteBus_req_bits_setIdx,
  input  [18:0] io_metaWriteBus_req_bits_data_tag,
  input         io_metaWriteBus_req_bits_data_dirty,
  input  [3:0]  io_metaWriteBus_req_bits_waymask,
  input         io_dataWriteBus_req_valid,
  input  [9:0]  io_dataWriteBus_req_bits_setIdx,
  input  [63:0] io_dataWriteBus_req_bits_data_data,
  input  [3:0]  io_dataWriteBus_req_bits_waymask,
  input         DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[Cache.scala 162:31]
  wire [6:0] addr_index = io_in_bits_req_addr[12:6]; // @[Cache.scala 162:31]
  wire [18:0] addr_tag = io_in_bits_req_addr[31:13]; // @[Cache.scala 162:31]
  wire  _T_5 = io_in_valid & io_metaWriteBus_req_valid; // @[Cache.scala 164:35]
  wire  _T_12 = io_metaWriteBus_req_bits_setIdx == addr_index; // @[Cache.scala 164:99]
  wire  isForwardMeta = _T_5 & _T_12; // @[Cache.scala 164:64]
  reg  isForwardMetaReg; // @[Cache.scala 165:33]
  wire  _GEN_0 = isForwardMeta | isForwardMetaReg; // @[Cache.scala 166:24]
  wire  _T_13 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire  _T_14 = ~io_in_valid; // @[Cache.scala 167:25]
  wire  _T_15 = _T_13 | _T_14; // @[Cache.scala 167:22]
  reg [18:0] forwardMetaReg_data_tag; // @[Reg.scala 15:16]
  reg  forwardMetaReg_data_dirty; // @[Reg.scala 15:16]
  reg [3:0] forwardMetaReg_waymask; // @[Reg.scala 15:16]
  wire [3:0] _GEN_2 = isForwardMeta ? io_metaWriteBus_req_bits_waymask : forwardMetaReg_waymask; // @[Reg.scala 16:19]
  wire  _GEN_3 = isForwardMeta ? io_metaWriteBus_req_bits_data_dirty : forwardMetaReg_data_dirty; // @[Reg.scala 16:19]
  wire [18:0] _GEN_5 = isForwardMeta ? io_metaWriteBus_req_bits_data_tag : forwardMetaReg_data_tag; // @[Reg.scala 16:19]
  wire  pickForwardMeta = isForwardMetaReg | isForwardMeta; // @[Cache.scala 171:42]
  wire  forwardWaymask_0 = _GEN_2[0]; // @[Cache.scala 173:61]
  wire  forwardWaymask_1 = _GEN_2[1]; // @[Cache.scala 173:61]
  wire  forwardWaymask_2 = _GEN_2[2]; // @[Cache.scala 173:61]
  wire  forwardWaymask_3 = _GEN_2[3]; // @[Cache.scala 173:61]
  wire  _T_16 = pickForwardMeta & forwardWaymask_0; // @[Cache.scala 175:39]
  wire [18:0] metaWay_0_tag = _T_16 ? _GEN_5 : io_metaReadResp_0_tag; // @[Cache.scala 175:22]
  wire  metaWay_0_valid = _T_16 | io_metaReadResp_0_valid; // @[Cache.scala 175:22]
  wire  _T_18 = pickForwardMeta & forwardWaymask_1; // @[Cache.scala 175:39]
  wire [18:0] metaWay_1_tag = _T_18 ? _GEN_5 : io_metaReadResp_1_tag; // @[Cache.scala 175:22]
  wire  metaWay_1_valid = _T_18 | io_metaReadResp_1_valid; // @[Cache.scala 175:22]
  wire  _T_20 = pickForwardMeta & forwardWaymask_2; // @[Cache.scala 175:39]
  wire [18:0] metaWay_2_tag = _T_20 ? _GEN_5 : io_metaReadResp_2_tag; // @[Cache.scala 175:22]
  wire  metaWay_2_valid = _T_20 | io_metaReadResp_2_valid; // @[Cache.scala 175:22]
  wire  _T_22 = pickForwardMeta & forwardWaymask_3; // @[Cache.scala 175:39]
  wire [18:0] metaWay_3_tag = _T_22 ? _GEN_5 : io_metaReadResp_3_tag; // @[Cache.scala 175:22]
  wire  metaWay_3_valid = _T_22 | io_metaReadResp_3_valid; // @[Cache.scala 175:22]
  wire  _T_24 = metaWay_0_tag == addr_tag; // @[Cache.scala 178:59]
  wire  _T_25 = metaWay_0_valid & _T_24; // @[Cache.scala 178:49]
  wire  _T_26 = _T_25 & io_in_valid; // @[Cache.scala 178:73]
  wire  _T_27 = metaWay_1_tag == addr_tag; // @[Cache.scala 178:59]
  wire  _T_28 = metaWay_1_valid & _T_27; // @[Cache.scala 178:49]
  wire  _T_29 = _T_28 & io_in_valid; // @[Cache.scala 178:73]
  wire  _T_30 = metaWay_2_tag == addr_tag; // @[Cache.scala 178:59]
  wire  _T_31 = metaWay_2_valid & _T_30; // @[Cache.scala 178:49]
  wire  _T_32 = _T_31 & io_in_valid; // @[Cache.scala 178:73]
  wire  _T_33 = metaWay_3_tag == addr_tag; // @[Cache.scala 178:59]
  wire  _T_34 = metaWay_3_valid & _T_33; // @[Cache.scala 178:49]
  wire  _T_35 = _T_34 & io_in_valid; // @[Cache.scala 178:73]
  wire [3:0] hitVec = {_T_35,_T_32,_T_29,_T_26}; // @[Cache.scala 178:90]
  reg [63:0] _T_39; // @[LFSR64.scala 25:23]
  wire  _T_42 = _T_39[0] ^ _T_39[1]; // @[LFSR64.scala 26:23]
  wire  _T_44 = _T_42 ^ _T_39[3]; // @[LFSR64.scala 26:33]
  wire  _T_46 = _T_44 ^ _T_39[4]; // @[LFSR64.scala 26:43]
  wire  _T_47 = _T_39 == 64'h0; // @[LFSR64.scala 28:24]
  wire [63:0] _T_49 = {_T_46,_T_39[63:1]}; // @[Cat.scala 29:58]
  wire [3:0] victimWaymask = 4'h1 << _T_39[1:0]; // @[Cache.scala 179:42]
  wire  _T_52 = ~metaWay_0_valid; // @[Cache.scala 181:45]
  wire  _T_53 = ~metaWay_1_valid; // @[Cache.scala 181:45]
  wire  _T_54 = ~metaWay_2_valid; // @[Cache.scala 181:45]
  wire  _T_55 = ~metaWay_3_valid; // @[Cache.scala 181:45]
  wire [3:0] invalidVec = {_T_55,_T_54,_T_53,_T_52}; // @[Cache.scala 181:56]
  wire  hasInvalidWay = |invalidVec; // @[Cache.scala 182:34]
  wire  _T_59 = invalidVec >= 4'h8; // @[Cache.scala 183:45]
  wire  _T_60 = invalidVec >= 4'h4; // @[Cache.scala 184:20]
  wire  _T_61 = invalidVec >= 4'h2; // @[Cache.scala 185:20]
  wire [1:0] _T_62 = _T_61 ? 2'h2 : 2'h1; // @[Cache.scala 185:8]
  wire [2:0] _T_63 = _T_60 ? 3'h4 : {{1'd0}, _T_62}; // @[Cache.scala 184:8]
  wire [3:0] refillInvalidWaymask = _T_59 ? 4'h8 : {{1'd0}, _T_63}; // @[Cache.scala 183:33]
  wire [3:0] _T_64 = hasInvalidWay ? refillInvalidWaymask : victimWaymask; // @[Cache.scala 188:49]
  wire [3:0] waymask = io_out_bits_hit ? hitVec : _T_64; // @[Cache.scala 188:20]
  wire [1:0] _T_69 = waymask[0] + waymask[1]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_71 = waymask[2] + waymask[3]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_73 = _T_69 + _T_71; // @[Bitwise.scala 47:55]
  wire  _T_75 = _T_73 > 3'h1; // @[Cache.scala 189:26]
  reg [63:0] _T_76; // @[GTimer.scala 24:20]
  wire [63:0] _T_78 = _T_76 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_82 = ~reset; // @[Debug.scala 56:24]
  reg [63:0] _T_85; // @[GTimer.scala 24:20]
  wire [63:0] _T_87 = _T_85 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_94; // @[GTimer.scala 24:20]
  wire [63:0] _T_96 = _T_94 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_103; // @[GTimer.scala 24:20]
  wire [63:0] _T_105 = _T_103 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_112; // @[GTimer.scala 24:20]
  wire [63:0] _T_114 = _T_112 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_121; // @[GTimer.scala 24:20]
  wire [63:0] _T_123 = _T_121 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_130; // @[GTimer.scala 24:20]
  wire [63:0] _T_132 = _T_130 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_139; // @[GTimer.scala 24:20]
  wire [63:0] _T_141 = _T_139 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_148; // @[GTimer.scala 24:20]
  wire [63:0] _T_150 = _T_148 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_157; // @[GTimer.scala 24:20]
  wire [63:0] _T_159 = _T_157 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_177; // @[GTimer.scala 24:20]
  wire [63:0] _T_179 = _T_177 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_197 = io_in_valid & _T_75; // @[Cache.scala 196:24]
  wire  _T_198 = ~_T_197; // @[Cache.scala 196:10]
  wire  _T_200 = _T_198 | reset; // @[Cache.scala 196:9]
  wire  _T_201 = ~_T_200; // @[Cache.scala 196:9]
  wire  _T_202 = |hitVec; // @[Cache.scala 199:44]
  wire [31:0] _T_204 = io_in_bits_req_addr ^ 32'h30000000; // @[NutCore.scala 86:11]
  wire  _T_206 = _T_204[31:28] == 4'h0; // @[NutCore.scala 86:44]
  wire [31:0] _T_207 = io_in_bits_req_addr ^ 32'h40000000; // @[NutCore.scala 86:11]
  wire  _T_209 = _T_207[31:30] == 2'h0; // @[NutCore.scala 86:44]
  wire [9:0] _T_223 = {addr_index,addr_wordIndex}; // @[Cat.scala 29:58]
  wire  _T_224 = io_dataWriteBus_req_bits_setIdx == _T_223; // @[Cache.scala 205:30]
  wire  _T_225 = io_dataWriteBus_req_valid & _T_224; // @[Cache.scala 205:13]
  wire  isForwardData = io_in_valid & _T_225; // @[Cache.scala 204:35]
  reg  isForwardDataReg; // @[Cache.scala 207:33]
  wire  _GEN_8 = isForwardData | isForwardDataReg; // @[Cache.scala 208:24]
  reg [63:0] forwardDataReg_data_data; // @[Reg.scala 15:16]
  reg [3:0] forwardDataReg_waymask; // @[Reg.scala 15:16]
  wire  _T_232 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  reg [63:0] _T_235; // @[GTimer.scala 24:20]
  wire [63:0] _T_237 = _T_235 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_250; // @[GTimer.scala 24:20]
  wire [63:0] _T_252 = _T_250 + 64'h1; // @[GTimer.scala 25:12]
  wire  _GEN_13 = _T_75 & DISPLAY_ENABLE; // @[Debug.scala 56:24]
  assign io_in_ready = _T_14 | _T_232; // @[Cache.scala 216:15]
  assign io_out_valid = io_in_valid; // @[Cache.scala 215:16]
  assign io_out_bits_req_addr = io_in_bits_req_addr; // @[Cache.scala 214:19]
  assign io_out_bits_req_size = io_in_bits_req_size; // @[Cache.scala 214:19]
  assign io_out_bits_req_cmd = io_in_bits_req_cmd; // @[Cache.scala 214:19]
  assign io_out_bits_req_wmask = io_in_bits_req_wmask; // @[Cache.scala 214:19]
  assign io_out_bits_req_wdata = io_in_bits_req_wdata; // @[Cache.scala 214:19]
  assign io_out_bits_metas_0_tag = _T_16 ? _GEN_5 : io_metaReadResp_0_tag; // @[Cache.scala 198:21]
  assign io_out_bits_metas_0_valid = _T_16 | io_metaReadResp_0_valid; // @[Cache.scala 198:21]
  assign io_out_bits_metas_0_dirty = _T_16 ? _GEN_3 : io_metaReadResp_0_dirty; // @[Cache.scala 198:21]
  assign io_out_bits_metas_1_tag = _T_18 ? _GEN_5 : io_metaReadResp_1_tag; // @[Cache.scala 198:21]
  assign io_out_bits_metas_1_valid = _T_18 | io_metaReadResp_1_valid; // @[Cache.scala 198:21]
  assign io_out_bits_metas_1_dirty = _T_18 ? _GEN_3 : io_metaReadResp_1_dirty; // @[Cache.scala 198:21]
  assign io_out_bits_metas_2_tag = _T_20 ? _GEN_5 : io_metaReadResp_2_tag; // @[Cache.scala 198:21]
  assign io_out_bits_metas_2_valid = _T_20 | io_metaReadResp_2_valid; // @[Cache.scala 198:21]
  assign io_out_bits_metas_2_dirty = _T_20 ? _GEN_3 : io_metaReadResp_2_dirty; // @[Cache.scala 198:21]
  assign io_out_bits_metas_3_tag = _T_22 ? _GEN_5 : io_metaReadResp_3_tag; // @[Cache.scala 198:21]
  assign io_out_bits_metas_3_valid = _T_22 | io_metaReadResp_3_valid; // @[Cache.scala 198:21]
  assign io_out_bits_metas_3_dirty = _T_22 ? _GEN_3 : io_metaReadResp_3_dirty; // @[Cache.scala 198:21]
  assign io_out_bits_datas_0_data = io_dataReadResp_0_data; // @[Cache.scala 201:21]
  assign io_out_bits_datas_1_data = io_dataReadResp_1_data; // @[Cache.scala 201:21]
  assign io_out_bits_datas_2_data = io_dataReadResp_2_data; // @[Cache.scala 201:21]
  assign io_out_bits_datas_3_data = io_dataReadResp_3_data; // @[Cache.scala 201:21]
  assign io_out_bits_hit = io_in_valid & _T_202; // @[Cache.scala 199:19]
  assign io_out_bits_waymask = io_out_bits_hit ? hitVec : _T_64; // @[Cache.scala 200:23]
  assign io_out_bits_mmio = _T_206 | _T_209; // @[Cache.scala 202:20]
  assign io_out_bits_isForwardData = isForwardDataReg | isForwardData; // @[Cache.scala 211:29]
  assign io_out_bits_forwardData_data_data = isForwardData ? io_dataWriteBus_req_bits_data_data : forwardDataReg_data_data; // @[Cache.scala 212:27]
  assign io_out_bits_forwardData_waymask = isForwardData ? io_dataWriteBus_req_bits_waymask : forwardDataReg_waymask; // @[Cache.scala 212:27]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  isForwardMetaReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  forwardMetaReg_data_tag = _RAND_1[18:0];
  _RAND_2 = {1{`RANDOM}};
  forwardMetaReg_data_dirty = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  forwardMetaReg_waymask = _RAND_3[3:0];
  _RAND_4 = {2{`RANDOM}};
  _T_39 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  _T_76 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  _T_85 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  _T_94 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  _T_103 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  _T_112 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  _T_121 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  _T_130 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  _T_139 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  _T_148 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  _T_157 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  _T_177 = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  isForwardDataReg = _RAND_16[0:0];
  _RAND_17 = {2{`RANDOM}};
  forwardDataReg_data_data = _RAND_17[63:0];
  _RAND_18 = {1{`RANDOM}};
  forwardDataReg_waymask = _RAND_18[3:0];
  _RAND_19 = {2{`RANDOM}};
  _T_235 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  _T_250 = _RAND_20[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      isForwardMetaReg <= 1'h0;
    end else if (_T_15) begin
      isForwardMetaReg <= 1'h0;
    end else begin
      isForwardMetaReg <= _GEN_0;
    end
    if (isForwardMeta) begin
      forwardMetaReg_data_tag <= io_metaWriteBus_req_bits_data_tag;
    end
    if (isForwardMeta) begin
      forwardMetaReg_data_dirty <= io_metaWriteBus_req_bits_data_dirty;
    end
    if (isForwardMeta) begin
      forwardMetaReg_waymask <= io_metaWriteBus_req_bits_waymask;
    end
    if (reset) begin
      _T_39 <= 64'h1234567887654321;
    end else if (_T_47) begin
      _T_39 <= 64'h1;
    end else begin
      _T_39 <= _T_49;
    end
    if (reset) begin
      _T_76 <= 64'h0;
    end else begin
      _T_76 <= _T_78;
    end
    if (reset) begin
      _T_85 <= 64'h0;
    end else begin
      _T_85 <= _T_87;
    end
    if (reset) begin
      _T_94 <= 64'h0;
    end else begin
      _T_94 <= _T_96;
    end
    if (reset) begin
      _T_103 <= 64'h0;
    end else begin
      _T_103 <= _T_105;
    end
    if (reset) begin
      _T_112 <= 64'h0;
    end else begin
      _T_112 <= _T_114;
    end
    if (reset) begin
      _T_121 <= 64'h0;
    end else begin
      _T_121 <= _T_123;
    end
    if (reset) begin
      _T_130 <= 64'h0;
    end else begin
      _T_130 <= _T_132;
    end
    if (reset) begin
      _T_139 <= 64'h0;
    end else begin
      _T_139 <= _T_141;
    end
    if (reset) begin
      _T_148 <= 64'h0;
    end else begin
      _T_148 <= _T_150;
    end
    if (reset) begin
      _T_157 <= 64'h0;
    end else begin
      _T_157 <= _T_159;
    end
    if (reset) begin
      _T_177 <= 64'h0;
    end else begin
      _T_177 <= _T_179;
    end
    if (reset) begin
      isForwardDataReg <= 1'h0;
    end else if (_T_15) begin
      isForwardDataReg <= 1'h0;
    end else begin
      isForwardDataReg <= _GEN_8;
    end
    if (isForwardData) begin
      forwardDataReg_data_data <= io_dataWriteBus_req_bits_data_data;
    end
    if (isForwardData) begin
      forwardDataReg_waymask <= io_dataWriteBus_req_bits_waymask;
    end
    if (reset) begin
      _T_235 <= 64'h0;
    end else begin
      _T_235 <= _T_237;
    end
    if (reset) begin
      _T_250 <= 64'h0;
    end else begin
      _T_250 <= _T_252;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_1: ",_T_76); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] metaWay %x metat %x reqt %x\n",metaWay_0_valid,metaWay_0_tag,addr_tag); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_1: ",_T_85); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] metaWay %x metat %x reqt %x\n",metaWay_1_valid,metaWay_1_tag,addr_tag); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_1: ",_T_94); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] metaWay %x metat %x reqt %x\n",metaWay_2_valid,metaWay_2_tag,addr_tag); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_1: ",_T_103); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] metaWay %x metat %x reqt %x\n",metaWay_3_valid,metaWay_3_tag,addr_tag); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_1: ",_T_112); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] metaReadResp %x metat %x reqt %x\n",io_metaReadResp_0_valid,io_metaReadResp_0_tag,addr_tag); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_1: ",_T_121); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] metaReadResp %x metat %x reqt %x\n",io_metaReadResp_1_valid,io_metaReadResp_1_tag,addr_tag); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_1: ",_T_130); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] metaReadResp %x metat %x reqt %x\n",io_metaReadResp_2_valid,io_metaReadResp_2_tag,addr_tag); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_1: ",_T_139); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] metaReadResp %x metat %x reqt %x\n",io_metaReadResp_3_valid,io_metaReadResp_3_tag,addr_tag); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_1: ",_T_148); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] forwardMetaReg isForwardMetaReg %x %x metat %x wm %b\n",isForwardMetaReg,1'h1,forwardMetaReg_data_tag,forwardMetaReg_waymask); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_1: ",_T_157); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] forwardMeta isForwardMeta %x %x metat %x wm %b\n",isForwardMeta,1'h1,io_metaWriteBus_req_bits_data_tag,io_metaWriteBus_req_bits_waymask); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_1: ",_T_177); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] hit %b wmask %b hitvec %b\n",io_out_bits_hit,_GEN_2,hitVec); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_201) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Cache.scala:196 assert(!(io.in.valid && PopCount(waymask) > 1.U))\n"); // @[Cache.scala 196:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_201) begin
          $fatal; // @[Cache.scala 196:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_1: ",_T_235); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_82) begin
          $fwrite(32'h80000002,"[isFD:%d isFDreg:%d inFire:%d invalid:%d \n",isForwardData,isForwardDataReg,_T_13,io_in_valid); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_1: ",_T_250); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_82) begin
          $fwrite(32'h80000002,"[isFM:%d isFMreg:%d metawreq:%x widx:%x ridx:%x \n",isForwardMeta,isForwardMetaReg,io_metaWriteBus_req_valid,io_metaWriteBus_req_bits_setIdx,addr_index); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CacheStage3_1(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_req_addr,
  input  [2:0]  io_in_bits_req_size,
  input  [3:0]  io_in_bits_req_cmd,
  input  [7:0]  io_in_bits_req_wmask,
  input  [63:0] io_in_bits_req_wdata,
  input  [18:0] io_in_bits_metas_0_tag,
  input         io_in_bits_metas_0_valid,
  input         io_in_bits_metas_0_dirty,
  input  [18:0] io_in_bits_metas_1_tag,
  input         io_in_bits_metas_1_valid,
  input         io_in_bits_metas_1_dirty,
  input  [18:0] io_in_bits_metas_2_tag,
  input         io_in_bits_metas_2_valid,
  input         io_in_bits_metas_2_dirty,
  input  [18:0] io_in_bits_metas_3_tag,
  input         io_in_bits_metas_3_valid,
  input         io_in_bits_metas_3_dirty,
  input  [63:0] io_in_bits_datas_0_data,
  input  [63:0] io_in_bits_datas_1_data,
  input  [63:0] io_in_bits_datas_2_data,
  input  [63:0] io_in_bits_datas_3_data,
  input         io_in_bits_hit,
  input  [3:0]  io_in_bits_waymask,
  input         io_in_bits_mmio,
  input         io_in_bits_isForwardData,
  input  [63:0] io_in_bits_forwardData_data_data,
  input  [3:0]  io_in_bits_forwardData_waymask,
  input         io_out_ready,
  output        io_out_valid,
  output [3:0]  io_out_bits_cmd,
  output [63:0] io_out_bits_rdata,
  output        io_isFinish,
  input         io_dataReadBus_req_ready,
  output        io_dataReadBus_req_valid,
  output [9:0]  io_dataReadBus_req_bits_setIdx,
  input  [63:0] io_dataReadBus_resp_data_0_data,
  input  [63:0] io_dataReadBus_resp_data_1_data,
  input  [63:0] io_dataReadBus_resp_data_2_data,
  input  [63:0] io_dataReadBus_resp_data_3_data,
  output        io_dataWriteBus_req_valid,
  output [9:0]  io_dataWriteBus_req_bits_setIdx,
  output [63:0] io_dataWriteBus_req_bits_data_data,
  output [3:0]  io_dataWriteBus_req_bits_waymask,
  output        io_metaWriteBus_req_valid,
  output [6:0]  io_metaWriteBus_req_bits_setIdx,
  output [18:0] io_metaWriteBus_req_bits_data_tag,
  output        io_metaWriteBus_req_bits_data_valid,
  output        io_metaWriteBus_req_bits_data_dirty,
  output [3:0]  io_metaWriteBus_req_bits_waymask,
  input         io_mem_req_ready,
  output        io_mem_req_valid,
  output [31:0] io_mem_req_bits_addr,
  output [2:0]  io_mem_req_bits_size,
  output [3:0]  io_mem_req_bits_cmd,
  output [7:0]  io_mem_req_bits_wmask,
  output [63:0] io_mem_req_bits_wdata,
  output        io_mem_resp_ready,
  input         io_mem_resp_valid,
  input  [3:0]  io_mem_resp_bits_cmd,
  input  [63:0] io_mem_resp_bits_rdata,
  input         io_mmio_req_ready,
  output        io_mmio_req_valid,
  output [31:0] io_mmio_req_bits_addr,
  output [2:0]  io_mmio_req_bits_size,
  output [3:0]  io_mmio_req_bits_cmd,
  output [7:0]  io_mmio_req_bits_wmask,
  output [63:0] io_mmio_req_bits_wdata,
  output        io_mmio_resp_ready,
  input         io_mmio_resp_valid,
  input  [63:0] io_mmio_resp_bits_rdata,
  output        io_cohResp_valid,
  output [3:0]  io_cohResp_bits_cmd,
  output [63:0] io_cohResp_bits_rdata,
  output        io_dataReadRespToL1,
  output        mmio_0,
  input         DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
`endif // RANDOMIZE_REG_INIT
  wire  metaWriteArb_io_in_0_valid; // @[Cache.scala 241:28]
  wire [6:0] metaWriteArb_io_in_0_bits_setIdx; // @[Cache.scala 241:28]
  wire [18:0] metaWriteArb_io_in_0_bits_data_tag; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_in_0_bits_data_dirty; // @[Cache.scala 241:28]
  wire [3:0] metaWriteArb_io_in_0_bits_waymask; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_in_1_valid; // @[Cache.scala 241:28]
  wire [6:0] metaWriteArb_io_in_1_bits_setIdx; // @[Cache.scala 241:28]
  wire [18:0] metaWriteArb_io_in_1_bits_data_tag; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_in_1_bits_data_dirty; // @[Cache.scala 241:28]
  wire [3:0] metaWriteArb_io_in_1_bits_waymask; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_out_valid; // @[Cache.scala 241:28]
  wire [6:0] metaWriteArb_io_out_bits_setIdx; // @[Cache.scala 241:28]
  wire [18:0] metaWriteArb_io_out_bits_data_tag; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_out_bits_data_dirty; // @[Cache.scala 241:28]
  wire [3:0] metaWriteArb_io_out_bits_waymask; // @[Cache.scala 241:28]
  wire  dataWriteArb_io_in_0_valid; // @[Cache.scala 242:28]
  wire [9:0] dataWriteArb_io_in_0_bits_setIdx; // @[Cache.scala 242:28]
  wire [63:0] dataWriteArb_io_in_0_bits_data_data; // @[Cache.scala 242:28]
  wire [3:0] dataWriteArb_io_in_0_bits_waymask; // @[Cache.scala 242:28]
  wire  dataWriteArb_io_in_1_valid; // @[Cache.scala 242:28]
  wire [9:0] dataWriteArb_io_in_1_bits_setIdx; // @[Cache.scala 242:28]
  wire [63:0] dataWriteArb_io_in_1_bits_data_data; // @[Cache.scala 242:28]
  wire [3:0] dataWriteArb_io_in_1_bits_waymask; // @[Cache.scala 242:28]
  wire  dataWriteArb_io_out_valid; // @[Cache.scala 242:28]
  wire [9:0] dataWriteArb_io_out_bits_setIdx; // @[Cache.scala 242:28]
  wire [63:0] dataWriteArb_io_out_bits_data_data; // @[Cache.scala 242:28]
  wire [3:0] dataWriteArb_io_out_bits_waymask; // @[Cache.scala 242:28]
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[Cache.scala 245:31]
  wire [6:0] addr_index = io_in_bits_req_addr[12:6]; // @[Cache.scala 245:31]
  wire [18:0] addr_tag = io_in_bits_req_addr[31:13]; // @[Cache.scala 245:31]
  wire  mmio = io_in_valid & io_in_bits_mmio; // @[Cache.scala 246:26]
  wire  hit = io_in_valid & io_in_bits_hit; // @[Cache.scala 247:25]
  wire  _T_5 = ~io_in_bits_hit; // @[Cache.scala 248:29]
  wire  miss = io_in_valid & _T_5; // @[Cache.scala 248:26]
  wire  _T_7 = io_in_bits_req_cmd == 4'h8; // @[SimpleBus.scala 79:23]
  wire  probe = io_in_valid & _T_7; // @[Cache.scala 249:39]
  wire  _T_8 = io_in_bits_req_cmd == 4'h2; // @[SimpleBus.scala 76:27]
  wire  hitReadBurst = hit & _T_8; // @[Cache.scala 250:26]
  wire [20:0] _T_14 = {io_in_bits_metas_0_tag,io_in_bits_metas_0_valid,io_in_bits_metas_0_dirty}; // @[Mux.scala 27:72]
  wire [20:0] _T_15 = io_in_bits_waymask[0] ? _T_14 : 21'h0; // @[Mux.scala 27:72]
  wire [20:0] _T_17 = {io_in_bits_metas_1_tag,io_in_bits_metas_1_valid,io_in_bits_metas_1_dirty}; // @[Mux.scala 27:72]
  wire [20:0] _T_18 = io_in_bits_waymask[1] ? _T_17 : 21'h0; // @[Mux.scala 27:72]
  wire [20:0] _T_20 = {io_in_bits_metas_2_tag,io_in_bits_metas_2_valid,io_in_bits_metas_2_dirty}; // @[Mux.scala 27:72]
  wire [20:0] _T_21 = io_in_bits_waymask[2] ? _T_20 : 21'h0; // @[Mux.scala 27:72]
  wire [20:0] _T_23 = {io_in_bits_metas_3_tag,io_in_bits_metas_3_valid,io_in_bits_metas_3_dirty}; // @[Mux.scala 27:72]
  wire [20:0] _T_24 = io_in_bits_waymask[3] ? _T_23 : 21'h0; // @[Mux.scala 27:72]
  wire [20:0] _T_25 = _T_15 | _T_18; // @[Mux.scala 27:72]
  wire [20:0] _T_26 = _T_25 | _T_21; // @[Mux.scala 27:72]
  wire [20:0] _T_27 = _T_26 | _T_24; // @[Mux.scala 27:72]
  wire  meta_dirty = _T_27[0]; // @[Mux.scala 27:72]
  wire [18:0] meta_tag = _T_27[20:2]; // @[Mux.scala 27:72]
  wire  _T_32 = mmio & hit; // @[Cache.scala 252:17]
  wire  _T_33 = ~_T_32; // @[Cache.scala 252:10]
  wire  _T_35 = _T_33 | reset; // @[Cache.scala 252:9]
  wire  _T_36 = ~_T_35; // @[Cache.scala 252:9]
  wire  _T_37 = io_in_bits_waymask == io_in_bits_forwardData_waymask; // @[Cache.scala 260:71]
  wire  useForwardData = io_in_bits_isForwardData & _T_37; // @[Cache.scala 260:49]
  wire [63:0] _T_42 = io_in_bits_waymask[0] ? io_in_bits_datas_0_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_43 = io_in_bits_waymask[1] ? io_in_bits_datas_1_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_44 = io_in_bits_waymask[2] ? io_in_bits_datas_2_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_45 = io_in_bits_waymask[3] ? io_in_bits_datas_3_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_46 = _T_42 | _T_43; // @[Mux.scala 27:72]
  wire [63:0] _T_47 = _T_46 | _T_44; // @[Mux.scala 27:72]
  wire [63:0] _T_48 = _T_47 | _T_45; // @[Mux.scala 27:72]
  wire [63:0] dataRead = useForwardData ? io_in_bits_forwardData_data_data : _T_48; // @[Cache.scala 262:21]
  wire [7:0] _T_64 = io_in_bits_req_wmask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_66 = io_in_bits_req_wmask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_68 = io_in_bits_req_wmask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_70 = io_in_bits_req_wmask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_72 = io_in_bits_req_wmask[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_74 = io_in_bits_req_wmask[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_76 = io_in_bits_req_wmask[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_78 = io_in_bits_req_wmask[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_85 = {_T_78,_T_76,_T_74,_T_72,_T_70,_T_68,_T_66,_T_64}; // @[Cat.scala 29:58]
  wire [63:0] wordMask = io_in_bits_req_cmd[0] ? _T_85 : 64'h0; // @[Cache.scala 263:21]
  reg [2:0] value; // @[Counter.scala 29:33]
  wire  _T_86 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_87 = io_in_bits_req_cmd == 4'h3; // @[Cache.scala 266:34]
  wire  _T_88 = io_in_bits_req_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_89 = _T_87 | _T_88; // @[Cache.scala 266:62]
  wire  _T_90 = _T_86 & _T_89; // @[Cache.scala 266:22]
  wire [2:0] _T_93 = value + 3'h1; // @[Counter.scala 39:22]
  wire [2:0] _GEN_0 = _T_90 ? _T_93 : value; // @[Cache.scala 266:85]
  wire  hitWrite = hit & io_in_bits_req_cmd[0]; // @[Cache.scala 270:22]
  wire [63:0] _T_96 = io_in_bits_req_wdata & wordMask; // @[BitUtils.scala 32:13]
  wire [63:0] _T_97 = ~wordMask; // @[BitUtils.scala 32:38]
  wire [63:0] _T_98 = dataRead & _T_97; // @[BitUtils.scala 32:36]
  wire [63:0] dataHitWriteBus_req_bits_data_data = _T_96 | _T_98; // @[BitUtils.scala 32:25]
  wire [2:0] _T_103 = _T_89 ? value : addr_wordIndex; // @[Cache.scala 273:51]
  wire [9:0] dataHitWriteBus_req_bits_setIdx = {addr_index,_T_103}; // @[Cat.scala 29:58]
  wire  _T_105 = ~meta_dirty; // @[Cache.scala 276:25]
  wire  metaHitWriteBus_req_valid = hitWrite & _T_105; // @[Cache.scala 276:22]
  reg [3:0] state; // @[Cache.scala 281:22]
  reg [2:0] value_1; // @[Counter.scala 29:33]
  reg [2:0] value_2; // @[Counter.scala 29:33]
  reg [1:0] state2; // @[Cache.scala 291:23]
  wire  _T_118 = state == 4'h3; // @[Cache.scala 293:39]
  wire  _T_119 = state == 4'h8; // @[Cache.scala 293:66]
  wire  _T_120 = _T_118 | _T_119; // @[Cache.scala 293:57]
  wire  _T_121 = state2 == 2'h0; // @[Cache.scala 293:92]
  wire [2:0] _T_124 = _T_119 ? value_1 : value_2; // @[Cache.scala 294:33]
  wire  _T_126 = state2 == 2'h1; // @[Cache.scala 295:60]
  reg [63:0] dataWay_0_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_1_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_2_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_3_data; // @[Reg.scala 15:16]
  wire [63:0] _T_131 = io_in_bits_waymask[0] ? dataWay_0_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_132 = io_in_bits_waymask[1] ? dataWay_1_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_133 = io_in_bits_waymask[2] ? dataWay_2_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_134 = io_in_bits_waymask[3] ? dataWay_3_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_135 = _T_131 | _T_132; // @[Mux.scala 27:72]
  wire [63:0] _T_136 = _T_135 | _T_133; // @[Mux.scala 27:72]
  wire  _T_141 = 2'h0 == state2; // @[Conditional.scala 37:30]
  wire  _T_142 = io_dataReadBus_req_ready & io_dataReadBus_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_143 = 2'h1 == state2; // @[Conditional.scala 37:30]
  wire  _T_144 = 2'h2 == state2; // @[Conditional.scala 37:30]
  wire  _T_145 = io_mem_req_ready & io_mem_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_147 = _T_145 | io_cohResp_valid; // @[Cache.scala 301:46]
  wire  _T_148 = hitReadBurst & io_out_ready; // @[Cache.scala 301:83]
  wire  _T_149 = _T_147 | _T_148; // @[Cache.scala 301:67]
  wire [31:0] raddr = {io_in_bits_req_addr[31:3],3'h0}; // @[Cat.scala 29:58]
  wire [31:0] waddr = {meta_tag,addr_index,6'h0}; // @[Cat.scala 29:58]
  wire  _T_152 = state == 4'h1; // @[Cache.scala 309:23]
  wire  _T_153 = value_2 == 3'h7; // @[Cache.scala 310:29]
  wire [2:0] _T_154 = _T_153 ? 3'h7 : 3'h3; // @[Cache.scala 310:8]
  wire [2:0] cmd = _T_152 ? 3'h2 : _T_154; // @[Cache.scala 309:16]
  wire  _T_160 = state2 == 2'h2; // @[Cache.scala 316:89]
  wire  _T_161 = _T_118 & _T_160; // @[Cache.scala 316:78]
  reg  afterFirstRead; // @[Cache.scala 323:31]
  reg  alreadyOutFire; // @[Reg.scala 27:20]
  wire  _GEN_12 = _T_86 | alreadyOutFire; // @[Reg.scala 28:19]
  wire  _T_165 = ~afterFirstRead; // @[Cache.scala 325:22]
  wire  _T_166 = io_mem_resp_ready & io_mem_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_167 = _T_165 & _T_166; // @[Cache.scala 325:38]
  wire  _T_168 = state == 4'h2; // @[Cache.scala 325:70]
  wire  readingFirst = _T_167 & _T_168; // @[Cache.scala 325:60]
  wire  _T_170 = state == 4'h6; // @[Cache.scala 327:52]
  wire  _T_171 = mmio ? _T_170 : readingFirst; // @[Cache.scala 327:39]
  reg [63:0] inRdataRegDemand; // @[Reg.scala 15:16]
  wire  _T_172 = state == 4'h0; // @[Cache.scala 330:31]
  wire  _T_173 = _T_172 & probe; // @[Cache.scala 330:43]
  wire  _T_176 = _T_119 & _T_160; // @[Cache.scala 331:46]
  wire  _T_180 = _T_119 & io_cohResp_valid; // @[Cache.scala 333:49]
  reg [2:0] _T_181; // @[Counter.scala 29:33]
  wire  _T_182 = _T_181 == 3'h7; // @[Counter.scala 38:24]
  wire [2:0] _T_184 = _T_181 + 3'h1; // @[Counter.scala 39:22]
  wire  releaseLast = _T_180 & _T_182; // @[Counter.scala 67:17]
  wire [2:0] _T_186 = releaseLast ? 3'h6 : 3'h0; // @[Cache.scala 334:54]
  wire [3:0] _T_187 = hit ? 4'hc : 4'h8; // @[Cache.scala 335:8]
  wire  respToL1Fire = _T_148 & _T_160; // @[Cache.scala 337:51]
  wire  _T_195 = _T_172 | _T_176; // @[Cache.scala 338:48]
  wire  _T_196 = _T_195 & hitReadBurst; // @[Cache.scala 338:96]
  wire  _T_197 = _T_196 & io_out_ready; // @[Cache.scala 338:112]
  reg [2:0] _T_198; // @[Counter.scala 29:33]
  wire  _T_199 = _T_198 == 3'h7; // @[Counter.scala 38:24]
  wire [2:0] _T_201 = _T_198 + 3'h1; // @[Counter.scala 39:22]
  wire  respToL1Last = _T_197 & _T_199; // @[Counter.scala 67:17]
  wire  _T_202 = 4'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_206 = addr_wordIndex == 3'h7; // @[Cache.scala 352:49]
  wire [2:0] _T_208 = addr_wordIndex + 3'h1; // @[Cache.scala 352:93]
  wire  _T_210 = miss | mmio; // @[Cache.scala 353:26]
  wire  _T_217 = 4'h5 == state; // @[Conditional.scala 37:30]
  wire  _T_218 = io_mmio_req_ready & io_mmio_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_219 = 4'h6 == state; // @[Conditional.scala 37:30]
  wire  _T_220 = io_mmio_resp_ready & io_mmio_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_221 = 4'h8 == state; // @[Conditional.scala 37:30]
  wire  _T_223 = io_cohResp_valid | respToL1Fire; // @[Cache.scala 362:31]
  wire [2:0] _T_226 = value_1 + 3'h1; // @[Counter.scala 39:22]
  wire  _T_228 = probe & io_cohResp_valid; // @[Cache.scala 363:19]
  wire  _T_229 = _T_228 & releaseLast; // @[Cache.scala 363:40]
  wire  _T_230 = respToL1Fire & respToL1Last; // @[Cache.scala 363:71]
  wire  _T_231 = _T_229 | _T_230; // @[Cache.scala 363:55]
  wire  _T_232 = 4'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_234 = 4'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_240 = io_mem_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire  _GEN_33 = _T_166 | afterFirstRead; // @[Cache.scala 372:33]
  wire  _T_241 = 4'h3 == state; // @[Conditional.scala 37:30]
  wire [2:0] _T_245 = value_2 + 3'h1; // @[Counter.scala 39:22]
  wire  _T_246 = io_mem_req_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_248 = _T_246 & _T_145; // @[Cache.scala 382:43]
  wire  _T_249 = 4'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_251 = 4'h7 == state; // @[Conditional.scala 37:30]
  wire [63:0] _T_255 = readingFirst ? wordMask : 64'h0; // @[Cache.scala 389:67]
  wire [63:0] _T_256 = io_in_bits_req_wdata & _T_255; // @[BitUtils.scala 32:13]
  wire [63:0] _T_257 = ~_T_255; // @[BitUtils.scala 32:38]
  wire [63:0] _T_258 = io_mem_resp_bits_rdata & _T_257; // @[BitUtils.scala 32:36]
  wire  dataRefillWriteBus_req_valid = _T_168 & _T_166; // @[Cache.scala 391:39]
  wire  metaRefillWriteBus_req_valid = dataRefillWriteBus_req_valid & _T_240; // @[Cache.scala 399:61]
  wire  _T_281 = ~io_in_bits_req_cmd[0]; // @[SimpleBus.scala 73:18]
  wire  _T_283 = ~io_in_bits_req_cmd[3]; // @[SimpleBus.scala 73:29]
  wire  _T_284 = _T_281 & _T_283; // @[SimpleBus.scala 73:26]
  wire [2:0] _T_286 = io_in_bits_req_cmd[0] ? 3'h5 : 3'h0; // @[Cache.scala 427:79]
  wire [2:0] _T_288 = _T_284 ? 3'h6 : _T_286; // @[Cache.scala 427:27]
  wire  _T_293 = state == 4'h7; // @[Cache.scala 433:48]
  wire  _T_308 = io_in_bits_req_cmd[0] | mmio; // @[Cache.scala 434:60]
  wire  _T_310 = ~alreadyOutFire; // @[Cache.scala 434:110]
  wire  _T_311 = afterFirstRead & _T_310; // @[Cache.scala 434:107]
  wire  _T_312 = _T_308 ? _T_293 : _T_311; // @[Cache.scala 434:45]
  wire  _T_313 = hit | _T_312; // @[Cache.scala 434:28]
  wire  _T_314 = probe ? 1'h0 : _T_313; // @[Cache.scala 434:8]
  wire  _T_320 = _T_119 & releaseLast; // @[Cache.scala 441:100]
  wire  _T_321 = miss ? _T_172 : _T_320; // @[Cache.scala 441:53]
  wire  _T_322 = io_cohResp_valid & _T_321; // @[Cache.scala 441:47]
  wire  _T_324 = hit | io_in_bits_req_cmd[0]; // @[Cache.scala 442:13]
  wire  _T_329 = _T_293 & _GEN_12; // @[Cache.scala 442:70]
  wire  _T_330 = _T_324 ? _T_86 : _T_329; // @[Cache.scala 442:8]
  wire  _T_333 = ~hitReadBurst; // @[Cache.scala 445:55]
  wire  _T_334 = _T_172 & _T_333; // @[Cache.scala 445:52]
  wire  _T_335 = io_out_ready & _T_334; // @[Cache.scala 445:31]
  wire  _T_336 = ~miss; // @[Cache.scala 445:73]
  wire  _T_337 = _T_335 & _T_336; // @[Cache.scala 445:70]
  wire  _T_338 = ~probe; // @[Cache.scala 445:82]
  wire  _T_341 = _T_172 & io_out_ready; // @[Cache.scala 446:60]
  wire  _T_345 = _T_341 | _T_176; // @[Cache.scala 446:76]
  wire  _T_347 = metaHitWriteBus_req_valid & metaRefillWriteBus_req_valid; // @[Cache.scala 448:38]
  wire  _T_348 = ~_T_347; // @[Cache.scala 448:10]
  wire  _T_350 = _T_348 | reset; // @[Cache.scala 448:9]
  wire  _T_351 = ~_T_350; // @[Cache.scala 448:9]
  wire  _T_352 = hitWrite & dataRefillWriteBus_req_valid; // @[Cache.scala 449:38]
  wire  _T_353 = ~_T_352; // @[Cache.scala 449:10]
  wire  _T_355 = _T_353 | reset; // @[Cache.scala 449:9]
  wire  _T_356 = ~_T_355; // @[Cache.scala 449:9]
  wire [255:0] _T_371 = {io_in_bits_datas_3_data,io_in_bits_datas_2_data,io_in_bits_datas_1_data,io_in_bits_datas_0_data}; // @[Cache.scala 451:465]
  reg [63:0] _T_372; // @[GTimer.scala 24:20]
  wire [63:0] _T_374 = _T_372 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_378 = ~reset; // @[Debug.scala 56:24]
  reg [63:0] _T_382; // @[GTimer.scala 24:20]
  wire [63:0] _T_384 = _T_382 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_385; // @[GTimer.scala 24:20]
  wire [63:0] _T_387 = _T_385 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_389 = io_metaWriteBus_req_valid & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  reg [63:0] _T_394; // @[GTimer.scala 24:20]
  wire [63:0] _T_396 = _T_394 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_403; // @[GTimer.scala 24:20]
  wire [63:0] _T_405 = _T_403 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_412; // @[GTimer.scala 24:20]
  wire [63:0] _T_414 = _T_412 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_424; // @[GTimer.scala 24:20]
  wire [63:0] _T_426 = _T_424 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_433; // @[GTimer.scala 24:20]
  wire [63:0] _T_435 = _T_433 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_443; // @[GTimer.scala 24:20]
  wire [63:0] _T_445 = _T_443 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_447 = io_dataWriteBus_req_valid & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  wire  _T_454 = _T_118 & _T_145; // @[Cache.scala 460:35]
  reg [63:0] _T_461; // @[GTimer.scala 24:20]
  wire [63:0] _T_463 = _T_461 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_465 = _T_454 & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  wire  _T_472 = _T_152 & _T_145; // @[Cache.scala 461:34]
  reg [63:0] _T_479; // @[GTimer.scala 24:20]
  wire [63:0] _T_481 = _T_479 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_483 = _T_472 & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  reg [63:0] _T_497; // @[GTimer.scala 24:20]
  wire [63:0] _T_499 = _T_497 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_501 = dataRefillWriteBus_req_valid & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  Arbiter metaWriteArb ( // @[Cache.scala 241:28]
    .io_in_0_valid(metaWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(metaWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_tag(metaWriteArb_io_in_0_bits_data_tag),
    .io_in_0_bits_data_dirty(metaWriteArb_io_in_0_bits_data_dirty),
    .io_in_0_bits_waymask(metaWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(metaWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(metaWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_tag(metaWriteArb_io_in_1_bits_data_tag),
    .io_in_1_bits_data_dirty(metaWriteArb_io_in_1_bits_data_dirty),
    .io_in_1_bits_waymask(metaWriteArb_io_in_1_bits_waymask),
    .io_out_valid(metaWriteArb_io_out_valid),
    .io_out_bits_setIdx(metaWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_tag(metaWriteArb_io_out_bits_data_tag),
    .io_out_bits_data_dirty(metaWriteArb_io_out_bits_data_dirty),
    .io_out_bits_waymask(metaWriteArb_io_out_bits_waymask)
  );
  Arbiter_1 dataWriteArb ( // @[Cache.scala 242:28]
    .io_in_0_valid(dataWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(dataWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_data(dataWriteArb_io_in_0_bits_data_data),
    .io_in_0_bits_waymask(dataWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(dataWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(dataWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_data(dataWriteArb_io_in_1_bits_data_data),
    .io_in_1_bits_waymask(dataWriteArb_io_in_1_bits_waymask),
    .io_out_valid(dataWriteArb_io_out_valid),
    .io_out_bits_setIdx(dataWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_data(dataWriteArb_io_out_bits_data_data),
    .io_out_bits_waymask(dataWriteArb_io_out_bits_waymask)
  );
  assign io_in_ready = _T_337 & _T_338; // @[Cache.scala 445:15]
  assign io_out_valid = io_in_valid & _T_314; // @[Cache.scala 432:16]
  assign io_out_bits_cmd = {{1'd0}, _T_288}; // @[Cache.scala 427:21]
  assign io_out_bits_rdata = hit ? dataRead : inRdataRegDemand; // @[Cache.scala 426:23]
  assign io_isFinish = probe ? _T_322 : _T_330; // @[Cache.scala 441:15]
  assign io_dataReadBus_req_valid = _T_120 & _T_121; // @[SRAMTemplate.scala 53:20]
  assign io_dataReadBus_req_bits_setIdx = {addr_index,_T_124}; // @[SRAMTemplate.scala 26:17]
  assign io_dataWriteBus_req_valid = dataWriteArb_io_out_valid; // @[Cache.scala 396:23]
  assign io_dataWriteBus_req_bits_setIdx = dataWriteArb_io_out_bits_setIdx; // @[Cache.scala 396:23]
  assign io_dataWriteBus_req_bits_data_data = dataWriteArb_io_out_bits_data_data; // @[Cache.scala 396:23]
  assign io_dataWriteBus_req_bits_waymask = dataWriteArb_io_out_bits_waymask; // @[Cache.scala 396:23]
  assign io_metaWriteBus_req_valid = metaWriteArb_io_out_valid; // @[Cache.scala 406:23]
  assign io_metaWriteBus_req_bits_setIdx = metaWriteArb_io_out_bits_setIdx; // @[Cache.scala 406:23]
  assign io_metaWriteBus_req_bits_data_tag = metaWriteArb_io_out_bits_data_tag; // @[Cache.scala 406:23]
  assign io_metaWriteBus_req_bits_data_valid = 1'h1; // @[Cache.scala 406:23]
  assign io_metaWriteBus_req_bits_data_dirty = metaWriteArb_io_out_bits_data_dirty; // @[Cache.scala 406:23]
  assign io_metaWriteBus_req_bits_waymask = metaWriteArb_io_out_bits_waymask; // @[Cache.scala 406:23]
  assign io_mem_req_valid = _T_152 | _T_161; // @[Cache.scala 316:20]
  assign io_mem_req_bits_addr = _T_152 ? raddr : waddr; // @[SimpleBus.scala 64:15]
  assign io_mem_req_bits_size = 3'h3; // @[SimpleBus.scala 66:15]
  assign io_mem_req_bits_cmd = {{1'd0}, cmd}; // @[SimpleBus.scala 65:14]
  assign io_mem_req_bits_wmask = 8'hff; // @[SimpleBus.scala 68:16]
  assign io_mem_req_bits_wdata = _T_136 | _T_134; // @[SimpleBus.scala 67:16]
  assign io_mem_resp_ready = 1'h1; // @[Cache.scala 315:21]
  assign io_mmio_req_valid = state == 4'h5; // @[Cache.scala 321:21]
  assign io_mmio_req_bits_addr = io_in_bits_req_addr; // @[Cache.scala 319:20]
  assign io_mmio_req_bits_size = io_in_bits_req_size; // @[Cache.scala 319:20]
  assign io_mmio_req_bits_cmd = io_in_bits_req_cmd; // @[Cache.scala 319:20]
  assign io_mmio_req_bits_wmask = io_in_bits_req_wmask; // @[Cache.scala 319:20]
  assign io_mmio_req_bits_wdata = io_in_bits_req_wdata; // @[Cache.scala 319:20]
  assign io_mmio_resp_ready = 1'h1; // @[Cache.scala 320:22]
  assign io_cohResp_valid = _T_173 | _T_176; // @[Cache.scala 330:20]
  assign io_cohResp_bits_cmd = _T_119 ? {{1'd0}, _T_186} : _T_187; // @[Cache.scala 334:23]
  assign io_cohResp_bits_rdata = _T_136 | _T_134; // @[Cache.scala 332:25]
  assign io_dataReadRespToL1 = hitReadBurst & _T_345; // @[Cache.scala 446:23]
  assign mmio_0 = mmio;
  assign metaWriteArb_io_in_0_valid = hitWrite & _T_105; // @[Cache.scala 404:25]
  assign metaWriteArb_io_in_0_bits_setIdx = io_in_bits_req_addr[12:6]; // @[Cache.scala 404:25]
  assign metaWriteArb_io_in_0_bits_data_tag = _T_27[20:2]; // @[Cache.scala 404:25]
  assign metaWriteArb_io_in_0_bits_data_dirty = 1'h1; // @[Cache.scala 404:25]
  assign metaWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[Cache.scala 404:25]
  assign metaWriteArb_io_in_1_valid = dataRefillWriteBus_req_valid & _T_240; // @[Cache.scala 405:25]
  assign metaWriteArb_io_in_1_bits_setIdx = io_in_bits_req_addr[12:6]; // @[Cache.scala 405:25]
  assign metaWriteArb_io_in_1_bits_data_tag = io_in_bits_req_addr[31:13]; // @[Cache.scala 405:25]
  assign metaWriteArb_io_in_1_bits_data_dirty = io_in_bits_req_cmd[0]; // @[Cache.scala 405:25]
  assign metaWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[Cache.scala 405:25]
  assign dataWriteArb_io_in_0_valid = hit & io_in_bits_req_cmd[0]; // @[Cache.scala 394:25]
  assign dataWriteArb_io_in_0_bits_setIdx = {addr_index,_T_103}; // @[Cache.scala 394:25]
  assign dataWriteArb_io_in_0_bits_data_data = _T_96 | _T_98; // @[Cache.scala 394:25]
  assign dataWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[Cache.scala 394:25]
  assign dataWriteArb_io_in_1_valid = _T_168 & _T_166; // @[Cache.scala 395:25]
  assign dataWriteArb_io_in_1_bits_setIdx = {addr_index,value_1}; // @[Cache.scala 395:25]
  assign dataWriteArb_io_in_1_bits_data_data = _T_256 | _T_258; // @[Cache.scala 395:25]
  assign dataWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[Cache.scala 395:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  value_2 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  state2 = _RAND_4[1:0];
  _RAND_5 = {2{`RANDOM}};
  dataWay_0_data = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  dataWay_1_data = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  dataWay_2_data = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  dataWay_3_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  afterFirstRead = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  alreadyOutFire = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  inRdataRegDemand = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  _T_181 = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  _T_198 = _RAND_13[2:0];
  _RAND_14 = {2{`RANDOM}};
  _T_372 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  _T_382 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  _T_385 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  _T_394 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  _T_403 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  _T_412 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  _T_424 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  _T_433 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  _T_443 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  _T_461 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  _T_479 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  _T_497 = _RAND_25[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 3'h0;
    end else if (_T_202) begin
      if (_T_90) begin
        value <= _T_93;
      end
    end else if (_T_217) begin
      if (_T_90) begin
        value <= _T_93;
      end
    end else if (_T_219) begin
      if (_T_90) begin
        value <= _T_93;
      end
    end else if (_T_221) begin
      if (_T_90) begin
        value <= _T_93;
      end
    end else if (_T_232) begin
      value <= _GEN_0;
    end else if (_T_234) begin
      if (_T_166) begin
        if (_T_87) begin
          value <= 3'h0;
        end else begin
          value <= _GEN_0;
        end
      end else begin
        value <= _GEN_0;
      end
    end else begin
      value <= _GEN_0;
    end
    if (reset) begin
      state <= 4'h0;
    end else if (_T_202) begin
      if (probe) begin
        if (io_cohResp_valid) begin
          if (hit) begin
            state <= 4'h8;
          end else begin
            state <= 4'h0;
          end
        end
      end else if (_T_148) begin
        state <= 4'h8;
      end else if (_T_210) begin
        if (mmio) begin
          state <= 4'h5;
        end else if (meta_dirty) begin
          state <= 4'h3;
        end else begin
          state <= 4'h1;
        end
      end
    end else if (_T_217) begin
      if (_T_218) begin
        state <= 4'h6;
      end
    end else if (_T_219) begin
      if (_T_220) begin
        state <= 4'h7;
      end
    end else if (_T_221) begin
      if (_T_231) begin
        state <= 4'h0;
      end
    end else if (_T_232) begin
      if (_T_145) begin
        state <= 4'h2;
      end
    end else if (_T_234) begin
      if (_T_166) begin
        if (_T_240) begin
          state <= 4'h7;
        end
      end
    end else if (_T_241) begin
      if (_T_248) begin
        state <= 4'h4;
      end
    end else if (_T_249) begin
      if (_T_166) begin
        state <= 4'h1;
      end
    end else if (_T_251) begin
      if (_GEN_12) begin
        state <= 4'h0;
      end
    end
    if (reset) begin
      value_1 <= 3'h0;
    end else if (_T_202) begin
      if (probe) begin
        if (io_cohResp_valid) begin
          value_1 <= addr_wordIndex;
        end
      end else if (_T_148) begin
        if (_T_206) begin
          value_1 <= 3'h0;
        end else begin
          value_1 <= _T_208;
        end
      end
    end else if (!(_T_217)) begin
      if (!(_T_219)) begin
        if (_T_221) begin
          if (_T_223) begin
            value_1 <= _T_226;
          end
        end else if (_T_232) begin
          if (_T_145) begin
            value_1 <= addr_wordIndex;
          end
        end else if (_T_234) begin
          if (_T_166) begin
            value_1 <= _T_226;
          end
        end
      end
    end
    if (reset) begin
      value_2 <= 3'h0;
    end else if (!(_T_202)) begin
      if (!(_T_217)) begin
        if (!(_T_219)) begin
          if (!(_T_221)) begin
            if (!(_T_232)) begin
              if (!(_T_234)) begin
                if (_T_241) begin
                  if (_T_145) begin
                    value_2 <= _T_245;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      state2 <= 2'h0;
    end else if (_T_141) begin
      if (_T_142) begin
        state2 <= 2'h1;
      end
    end else if (_T_143) begin
      state2 <= 2'h2;
    end else if (_T_144) begin
      if (_T_149) begin
        state2 <= 2'h0;
      end
    end
    if (_T_126) begin
      dataWay_0_data <= io_dataReadBus_resp_data_0_data;
    end
    if (_T_126) begin
      dataWay_1_data <= io_dataReadBus_resp_data_1_data;
    end
    if (_T_126) begin
      dataWay_2_data <= io_dataReadBus_resp_data_2_data;
    end
    if (_T_126) begin
      dataWay_3_data <= io_dataReadBus_resp_data_3_data;
    end
    if (reset) begin
      afterFirstRead <= 1'h0;
    end else if (_T_202) begin
      afterFirstRead <= 1'h0;
    end else if (!(_T_217)) begin
      if (!(_T_219)) begin
        if (!(_T_221)) begin
          if (!(_T_232)) begin
            if (_T_234) begin
              afterFirstRead <= _GEN_33;
            end
          end
        end
      end
    end
    if (reset) begin
      alreadyOutFire <= 1'h0;
    end else if (_T_202) begin
      alreadyOutFire <= 1'h0;
    end else begin
      alreadyOutFire <= _GEN_12;
    end
    if (_T_171) begin
      if (mmio) begin
        inRdataRegDemand <= io_mmio_resp_bits_rdata;
      end else begin
        inRdataRegDemand <= io_mem_resp_bits_rdata;
      end
    end
    if (reset) begin
      _T_181 <= 3'h0;
    end else if (_T_180) begin
      _T_181 <= _T_184;
    end
    if (reset) begin
      _T_198 <= 3'h0;
    end else if (_T_197) begin
      _T_198 <= _T_201;
    end
    if (reset) begin
      _T_372 <= 64'h0;
    end else begin
      _T_372 <= _T_374;
    end
    if (reset) begin
      _T_382 <= 64'h0;
    end else begin
      _T_382 <= _T_384;
    end
    if (reset) begin
      _T_385 <= 64'h0;
    end else begin
      _T_385 <= _T_387;
    end
    if (reset) begin
      _T_394 <= 64'h0;
    end else begin
      _T_394 <= _T_396;
    end
    if (reset) begin
      _T_403 <= 64'h0;
    end else begin
      _T_403 <= _T_405;
    end
    if (reset) begin
      _T_412 <= 64'h0;
    end else begin
      _T_412 <= _T_414;
    end
    if (reset) begin
      _T_424 <= 64'h0;
    end else begin
      _T_424 <= _T_426;
    end
    if (reset) begin
      _T_433 <= 64'h0;
    end else begin
      _T_433 <= _T_435;
    end
    if (reset) begin
      _T_443 <= 64'h0;
    end else begin
      _T_443 <= _T_445;
    end
    if (reset) begin
      _T_461 <= 64'h0;
    end else begin
      _T_461 <= _T_463;
    end
    if (reset) begin
      _T_479 <= 64'h0;
    end else begin
      _T_479 <= _T_481;
    end
    if (reset) begin
      _T_497 <= 64'h0;
    end else begin
      _T_497 <= _T_499;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_36) begin
          $fwrite(32'h80000002,"Assertion failed: MMIO request should not hit in cache\n    at Cache.scala:252 assert(!(mmio && hit), \"MMIO request should not hit in cache\")\n"); // @[Cache.scala 252:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_36) begin
          $fatal; // @[Cache.scala 252:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_351) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Cache.scala:448 assert(!(metaHitWriteBus.req.valid && metaRefillWriteBus.req.valid))\n"); // @[Cache.scala 448:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_351) begin
          $fatal; // @[Cache.scala 448:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_356) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Cache.scala:449 assert(!(dataHitWriteBus.req.valid && dataRefillWriteBus.req.valid))\n"); // @[Cache.scala 449:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_356) begin
          $fatal; // @[Cache.scala 449:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_378) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_1: ",_T_372); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_378) begin
          $fwrite(32'h80000002," metaread idx %x waymask %b metas %x%x:%x %x%x:%x %x%x:%x %x%x:%x %x\n",addr_index,io_in_bits_waymask,io_in_bits_metas_0_valid,io_in_bits_metas_0_dirty,io_in_bits_metas_0_tag,io_in_bits_metas_1_valid,io_in_bits_metas_1_dirty,io_in_bits_metas_1_tag,io_in_bits_metas_2_valid,io_in_bits_metas_2_dirty,io_in_bits_metas_2_tag,io_in_bits_metas_3_valid,io_in_bits_metas_3_dirty,io_in_bits_metas_3_tag,_T_371); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_389 & _T_378) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_1: ",_T_385); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_389 & _T_378) begin
          $fwrite(32'h80000002,"%d: [dcache S3]: metawrite idx %x wmask %b meta %x%x:%x\n",_T_382,io_metaWriteBus_req_bits_setIdx,io_metaWriteBus_req_bits_waymask,io_metaWriteBus_req_bits_data_valid,io_metaWriteBus_req_bits_data_dirty,io_metaWriteBus_req_bits_data_tag); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_378) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_1: ",_T_394); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_378) begin
          $fwrite(32'h80000002," in.ready = %d, in.valid = %d, hit = %x, state = %d, addr = %x cmd:%d probe:%d isFinish:%d\n",io_in_ready,io_in_valid,hit,state,io_in_bits_req_addr,io_in_bits_req_cmd,probe,io_isFinish); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_378) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_1: ",_T_403); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_378) begin
          $fwrite(32'h80000002," out.valid:%d rdata:%x cmd:%d user:%x id:%x \n",io_out_valid,io_out_bits_rdata,io_out_bits_cmd,1'h0,1'h0); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_378) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_1: ",_T_412); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_378) begin
          $fwrite(32'h80000002," DHW: (%d, %d), data:%x setIdx:%x MHW:(%d, %d)\n",hitWrite,1'h1,dataHitWriteBus_req_bits_data_data,dataHitWriteBus_req_bits_setIdx,metaHitWriteBus_req_valid,1'h1); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_378) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_1: ",_T_424); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_378) begin
          $fwrite(32'h80000002," DreadCache: %x \n",_T_371); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_378) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_1: ",_T_433); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_378) begin
          $fwrite(32'h80000002," useFD:%d isFD:%d FD:%x DreadArray:%x dataRead:%x inwaymask:%x FDwaymask:%x \n",useForwardData,io_in_bits_isForwardData,io_in_bits_forwardData_data_data,_T_48,dataRead,io_in_bits_waymask,io_in_bits_forwardData_waymask); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_447 & _T_378) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_1: ",_T_443); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_447 & _T_378) begin
          $fwrite(32'h80000002,"[WB] waymask: %b data:%x setIdx:%x\n",io_dataWriteBus_req_bits_waymask,io_dataWriteBus_req_bits_data_data,io_dataWriteBus_req_bits_setIdx); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_465 & _T_378) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_1: ",_T_461); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_465 & _T_378) begin
          $fwrite(32'h80000002,"[COUTW] cnt %x addr %x data %x cmd %x size %x wmask %x tag %x idx %x waymask %b \n",value_2,io_mem_req_bits_addr,io_mem_req_bits_wdata,io_mem_req_bits_cmd,io_mem_req_bits_size,io_mem_req_bits_wmask,addr_tag,addr_index,io_in_bits_waymask); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_483 & _T_378) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_1: ",_T_479); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_483 & _T_378) begin
          $fwrite(32'h80000002,"[COUTR] addr %x tag %x idx %x waymask %b \n",io_mem_req_bits_addr,addr_tag,addr_index,io_in_bits_waymask); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_501 & _T_378) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_1: ",_T_497); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_501 & _T_378) begin
          $fwrite(32'h80000002,"[COUTR] cnt %x data %x tag %x idx %x waymask %b \n",value_1,io_mem_resp_bits_rdata,addr_tag,addr_index,io_in_bits_waymask); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Arbiter_9(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input  [2:0]  io_in_0_bits_size,
  input  [3:0]  io_in_0_bits_cmd,
  input  [7:0]  io_in_0_bits_wmask,
  input  [63:0] io_in_0_bits_wdata,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input  [2:0]  io_in_1_bits_size,
  input  [3:0]  io_in_1_bits_cmd,
  input  [7:0]  io_in_1_bits_wmask,
  input  [63:0] io_in_1_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [2:0]  io_out_bits_size,
  output [3:0]  io_out_bits_cmd,
  output [7:0]  io_out_bits_wmask,
  output [63:0] io_out_bits_wdata
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  wire  _T_2 = ~grant_1; // @[Arbiter.scala 135:19]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:14]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_out_valid = _T_2 | io_in_1_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : io_in_1_bits_addr; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_size = io_in_0_valid ? io_in_0_bits_size : io_in_1_bits_size; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_cmd = io_in_0_valid ? io_in_0_bits_cmd : io_in_1_bits_cmd; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_wmask = io_in_0_valid ? io_in_0_bits_wmask : io_in_1_bits_wmask; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_wdata = io_in_0_valid ? io_in_0_bits_wdata : io_in_1_bits_wdata; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
endmodule
module Cache_1(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [2:0]  io_in_req_bits_size,
  input  [3:0]  io_in_req_bits_cmd,
  input  [7:0]  io_in_req_bits_wmask,
  input  [63:0] io_in_req_bits_wdata,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_mem_req_ready,
  output        io_out_mem_req_valid,
  output [31:0] io_out_mem_req_bits_addr,
  output [3:0]  io_out_mem_req_bits_cmd,
  output [63:0] io_out_mem_req_bits_wdata,
  input         io_out_mem_resp_valid,
  input  [3:0]  io_out_mem_resp_bits_cmd,
  input  [63:0] io_out_mem_resp_bits_rdata,
  output        io_out_coh_req_ready,
  input         io_out_coh_req_valid,
  input  [31:0] io_out_coh_req_bits_addr,
  input  [63:0] io_out_coh_req_bits_wdata,
  output        io_out_coh_resp_valid,
  output [3:0]  io_out_coh_resp_bits_cmd,
  output [63:0] io_out_coh_resp_bits_rdata,
  input         io_mmio_req_ready,
  output        io_mmio_req_valid,
  output [31:0] io_mmio_req_bits_addr,
  output [2:0]  io_mmio_req_bits_size,
  output [3:0]  io_mmio_req_bits_cmd,
  output [7:0]  io_mmio_req_bits_wmask,
  output [63:0] io_mmio_req_bits_wdata,
  input         io_mmio_resp_valid,
  input  [63:0] io_mmio_resp_bits_rdata,
  output        io_empty,
  output        mmio,
  input         DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
`endif // RANDOMIZE_REG_INIT
  wire  s1_clock; // @[Cache.scala 475:18]
  wire  s1_reset; // @[Cache.scala 475:18]
  wire  s1_io_in_ready; // @[Cache.scala 475:18]
  wire  s1_io_in_valid; // @[Cache.scala 475:18]
  wire [31:0] s1_io_in_bits_addr; // @[Cache.scala 475:18]
  wire [2:0] s1_io_in_bits_size; // @[Cache.scala 475:18]
  wire [3:0] s1_io_in_bits_cmd; // @[Cache.scala 475:18]
  wire [7:0] s1_io_in_bits_wmask; // @[Cache.scala 475:18]
  wire [63:0] s1_io_in_bits_wdata; // @[Cache.scala 475:18]
  wire  s1_io_out_ready; // @[Cache.scala 475:18]
  wire  s1_io_out_valid; // @[Cache.scala 475:18]
  wire [31:0] s1_io_out_bits_req_addr; // @[Cache.scala 475:18]
  wire [2:0] s1_io_out_bits_req_size; // @[Cache.scala 475:18]
  wire [3:0] s1_io_out_bits_req_cmd; // @[Cache.scala 475:18]
  wire [7:0] s1_io_out_bits_req_wmask; // @[Cache.scala 475:18]
  wire [63:0] s1_io_out_bits_req_wdata; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_req_ready; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_req_valid; // @[Cache.scala 475:18]
  wire [6:0] s1_io_metaReadBus_req_bits_setIdx; // @[Cache.scala 475:18]
  wire [18:0] s1_io_metaReadBus_resp_data_0_tag; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_0_valid; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_0_dirty; // @[Cache.scala 475:18]
  wire [18:0] s1_io_metaReadBus_resp_data_1_tag; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_1_valid; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_1_dirty; // @[Cache.scala 475:18]
  wire [18:0] s1_io_metaReadBus_resp_data_2_tag; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_2_valid; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_2_dirty; // @[Cache.scala 475:18]
  wire [18:0] s1_io_metaReadBus_resp_data_3_tag; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_3_valid; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_3_dirty; // @[Cache.scala 475:18]
  wire  s1_io_dataReadBus_req_ready; // @[Cache.scala 475:18]
  wire  s1_io_dataReadBus_req_valid; // @[Cache.scala 475:18]
  wire [9:0] s1_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 475:18]
  wire [63:0] s1_io_dataReadBus_resp_data_0_data; // @[Cache.scala 475:18]
  wire [63:0] s1_io_dataReadBus_resp_data_1_data; // @[Cache.scala 475:18]
  wire [63:0] s1_io_dataReadBus_resp_data_2_data; // @[Cache.scala 475:18]
  wire [63:0] s1_io_dataReadBus_resp_data_3_data; // @[Cache.scala 475:18]
  wire  s1_DISPLAY_ENABLE; // @[Cache.scala 475:18]
  wire  s2_clock; // @[Cache.scala 476:18]
  wire  s2_reset; // @[Cache.scala 476:18]
  wire  s2_io_in_ready; // @[Cache.scala 476:18]
  wire  s2_io_in_valid; // @[Cache.scala 476:18]
  wire [31:0] s2_io_in_bits_req_addr; // @[Cache.scala 476:18]
  wire [2:0] s2_io_in_bits_req_size; // @[Cache.scala 476:18]
  wire [3:0] s2_io_in_bits_req_cmd; // @[Cache.scala 476:18]
  wire [7:0] s2_io_in_bits_req_wmask; // @[Cache.scala 476:18]
  wire [63:0] s2_io_in_bits_req_wdata; // @[Cache.scala 476:18]
  wire  s2_io_out_ready; // @[Cache.scala 476:18]
  wire  s2_io_out_valid; // @[Cache.scala 476:18]
  wire [31:0] s2_io_out_bits_req_addr; // @[Cache.scala 476:18]
  wire [2:0] s2_io_out_bits_req_size; // @[Cache.scala 476:18]
  wire [3:0] s2_io_out_bits_req_cmd; // @[Cache.scala 476:18]
  wire [7:0] s2_io_out_bits_req_wmask; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_req_wdata; // @[Cache.scala 476:18]
  wire [18:0] s2_io_out_bits_metas_0_tag; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_0_valid; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_0_dirty; // @[Cache.scala 476:18]
  wire [18:0] s2_io_out_bits_metas_1_tag; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_1_valid; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_1_dirty; // @[Cache.scala 476:18]
  wire [18:0] s2_io_out_bits_metas_2_tag; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_2_valid; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_2_dirty; // @[Cache.scala 476:18]
  wire [18:0] s2_io_out_bits_metas_3_tag; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_3_valid; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_3_dirty; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_datas_0_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_datas_1_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_datas_2_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_datas_3_data; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_hit; // @[Cache.scala 476:18]
  wire [3:0] s2_io_out_bits_waymask; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_mmio; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_isForwardData; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_forwardData_data_data; // @[Cache.scala 476:18]
  wire [3:0] s2_io_out_bits_forwardData_waymask; // @[Cache.scala 476:18]
  wire [18:0] s2_io_metaReadResp_0_tag; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_0_valid; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_0_dirty; // @[Cache.scala 476:18]
  wire [18:0] s2_io_metaReadResp_1_tag; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_1_valid; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_1_dirty; // @[Cache.scala 476:18]
  wire [18:0] s2_io_metaReadResp_2_tag; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_2_valid; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_2_dirty; // @[Cache.scala 476:18]
  wire [18:0] s2_io_metaReadResp_3_tag; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_3_valid; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_3_dirty; // @[Cache.scala 476:18]
  wire [63:0] s2_io_dataReadResp_0_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_dataReadResp_1_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_dataReadResp_2_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_dataReadResp_3_data; // @[Cache.scala 476:18]
  wire  s2_io_metaWriteBus_req_valid; // @[Cache.scala 476:18]
  wire [6:0] s2_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 476:18]
  wire [18:0] s2_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 476:18]
  wire  s2_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 476:18]
  wire [3:0] s2_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 476:18]
  wire  s2_io_dataWriteBus_req_valid; // @[Cache.scala 476:18]
  wire [9:0] s2_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 476:18]
  wire [63:0] s2_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 476:18]
  wire [3:0] s2_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 476:18]
  wire  s2_DISPLAY_ENABLE; // @[Cache.scala 476:18]
  wire  s3_clock; // @[Cache.scala 477:18]
  wire  s3_reset; // @[Cache.scala 477:18]
  wire  s3_io_in_ready; // @[Cache.scala 477:18]
  wire  s3_io_in_valid; // @[Cache.scala 477:18]
  wire [31:0] s3_io_in_bits_req_addr; // @[Cache.scala 477:18]
  wire [2:0] s3_io_in_bits_req_size; // @[Cache.scala 477:18]
  wire [3:0] s3_io_in_bits_req_cmd; // @[Cache.scala 477:18]
  wire [7:0] s3_io_in_bits_req_wmask; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_req_wdata; // @[Cache.scala 477:18]
  wire [18:0] s3_io_in_bits_metas_0_tag; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_0_valid; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_0_dirty; // @[Cache.scala 477:18]
  wire [18:0] s3_io_in_bits_metas_1_tag; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_1_valid; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_1_dirty; // @[Cache.scala 477:18]
  wire [18:0] s3_io_in_bits_metas_2_tag; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_2_valid; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_2_dirty; // @[Cache.scala 477:18]
  wire [18:0] s3_io_in_bits_metas_3_tag; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_3_valid; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_3_dirty; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_datas_0_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_datas_1_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_datas_2_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_datas_3_data; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_hit; // @[Cache.scala 477:18]
  wire [3:0] s3_io_in_bits_waymask; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_mmio; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_isForwardData; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_forwardData_data_data; // @[Cache.scala 477:18]
  wire [3:0] s3_io_in_bits_forwardData_waymask; // @[Cache.scala 477:18]
  wire  s3_io_out_ready; // @[Cache.scala 477:18]
  wire  s3_io_out_valid; // @[Cache.scala 477:18]
  wire [3:0] s3_io_out_bits_cmd; // @[Cache.scala 477:18]
  wire [63:0] s3_io_out_bits_rdata; // @[Cache.scala 477:18]
  wire  s3_io_isFinish; // @[Cache.scala 477:18]
  wire  s3_io_dataReadBus_req_ready; // @[Cache.scala 477:18]
  wire  s3_io_dataReadBus_req_valid; // @[Cache.scala 477:18]
  wire [9:0] s3_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 477:18]
  wire [63:0] s3_io_dataReadBus_resp_data_0_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_dataReadBus_resp_data_1_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_dataReadBus_resp_data_2_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_dataReadBus_resp_data_3_data; // @[Cache.scala 477:18]
  wire  s3_io_dataWriteBus_req_valid; // @[Cache.scala 477:18]
  wire [9:0] s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 477:18]
  wire [63:0] s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 477:18]
  wire [3:0] s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 477:18]
  wire  s3_io_metaWriteBus_req_valid; // @[Cache.scala 477:18]
  wire [6:0] s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 477:18]
  wire [18:0] s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 477:18]
  wire  s3_io_metaWriteBus_req_bits_data_valid; // @[Cache.scala 477:18]
  wire  s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 477:18]
  wire [3:0] s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 477:18]
  wire  s3_io_mem_req_ready; // @[Cache.scala 477:18]
  wire  s3_io_mem_req_valid; // @[Cache.scala 477:18]
  wire [31:0] s3_io_mem_req_bits_addr; // @[Cache.scala 477:18]
  wire [2:0] s3_io_mem_req_bits_size; // @[Cache.scala 477:18]
  wire [3:0] s3_io_mem_req_bits_cmd; // @[Cache.scala 477:18]
  wire [7:0] s3_io_mem_req_bits_wmask; // @[Cache.scala 477:18]
  wire [63:0] s3_io_mem_req_bits_wdata; // @[Cache.scala 477:18]
  wire  s3_io_mem_resp_ready; // @[Cache.scala 477:18]
  wire  s3_io_mem_resp_valid; // @[Cache.scala 477:18]
  wire [3:0] s3_io_mem_resp_bits_cmd; // @[Cache.scala 477:18]
  wire [63:0] s3_io_mem_resp_bits_rdata; // @[Cache.scala 477:18]
  wire  s3_io_mmio_req_ready; // @[Cache.scala 477:18]
  wire  s3_io_mmio_req_valid; // @[Cache.scala 477:18]
  wire [31:0] s3_io_mmio_req_bits_addr; // @[Cache.scala 477:18]
  wire [2:0] s3_io_mmio_req_bits_size; // @[Cache.scala 477:18]
  wire [3:0] s3_io_mmio_req_bits_cmd; // @[Cache.scala 477:18]
  wire [7:0] s3_io_mmio_req_bits_wmask; // @[Cache.scala 477:18]
  wire [63:0] s3_io_mmio_req_bits_wdata; // @[Cache.scala 477:18]
  wire  s3_io_mmio_resp_ready; // @[Cache.scala 477:18]
  wire  s3_io_mmio_resp_valid; // @[Cache.scala 477:18]
  wire [63:0] s3_io_mmio_resp_bits_rdata; // @[Cache.scala 477:18]
  wire  s3_io_cohResp_valid; // @[Cache.scala 477:18]
  wire [3:0] s3_io_cohResp_bits_cmd; // @[Cache.scala 477:18]
  wire [63:0] s3_io_cohResp_bits_rdata; // @[Cache.scala 477:18]
  wire  s3_io_dataReadRespToL1; // @[Cache.scala 477:18]
  wire  s3_mmio_0; // @[Cache.scala 477:18]
  wire  s3_DISPLAY_ENABLE; // @[Cache.scala 477:18]
  wire  metaArray_clock; // @[Cache.scala 478:25]
  wire  metaArray_reset; // @[Cache.scala 478:25]
  wire  metaArray_io_r_0_req_ready; // @[Cache.scala 478:25]
  wire  metaArray_io_r_0_req_valid; // @[Cache.scala 478:25]
  wire [6:0] metaArray_io_r_0_req_bits_setIdx; // @[Cache.scala 478:25]
  wire [18:0] metaArray_io_r_0_resp_data_0_tag; // @[Cache.scala 478:25]
  wire  metaArray_io_r_0_resp_data_0_valid; // @[Cache.scala 478:25]
  wire  metaArray_io_r_0_resp_data_0_dirty; // @[Cache.scala 478:25]
  wire [18:0] metaArray_io_r_0_resp_data_1_tag; // @[Cache.scala 478:25]
  wire  metaArray_io_r_0_resp_data_1_valid; // @[Cache.scala 478:25]
  wire  metaArray_io_r_0_resp_data_1_dirty; // @[Cache.scala 478:25]
  wire [18:0] metaArray_io_r_0_resp_data_2_tag; // @[Cache.scala 478:25]
  wire  metaArray_io_r_0_resp_data_2_valid; // @[Cache.scala 478:25]
  wire  metaArray_io_r_0_resp_data_2_dirty; // @[Cache.scala 478:25]
  wire [18:0] metaArray_io_r_0_resp_data_3_tag; // @[Cache.scala 478:25]
  wire  metaArray_io_r_0_resp_data_3_valid; // @[Cache.scala 478:25]
  wire  metaArray_io_r_0_resp_data_3_dirty; // @[Cache.scala 478:25]
  wire  metaArray_io_w_req_valid; // @[Cache.scala 478:25]
  wire [6:0] metaArray_io_w_req_bits_setIdx; // @[Cache.scala 478:25]
  wire [18:0] metaArray_io_w_req_bits_data_tag; // @[Cache.scala 478:25]
  wire  metaArray_io_w_req_bits_data_dirty; // @[Cache.scala 478:25]
  wire [3:0] metaArray_io_w_req_bits_waymask; // @[Cache.scala 478:25]
  wire  dataArray_clock; // @[Cache.scala 479:25]
  wire  dataArray_reset; // @[Cache.scala 479:25]
  wire  dataArray_io_r_0_req_ready; // @[Cache.scala 479:25]
  wire  dataArray_io_r_0_req_valid; // @[Cache.scala 479:25]
  wire [9:0] dataArray_io_r_0_req_bits_setIdx; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r_0_resp_data_0_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r_0_resp_data_1_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r_0_resp_data_2_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r_0_resp_data_3_data; // @[Cache.scala 479:25]
  wire  dataArray_io_r_1_req_ready; // @[Cache.scala 479:25]
  wire  dataArray_io_r_1_req_valid; // @[Cache.scala 479:25]
  wire [9:0] dataArray_io_r_1_req_bits_setIdx; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r_1_resp_data_0_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r_1_resp_data_1_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r_1_resp_data_2_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r_1_resp_data_3_data; // @[Cache.scala 479:25]
  wire  dataArray_io_w_req_valid; // @[Cache.scala 479:25]
  wire [9:0] dataArray_io_w_req_bits_setIdx; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_w_req_bits_data_data; // @[Cache.scala 479:25]
  wire [3:0] dataArray_io_w_req_bits_waymask; // @[Cache.scala 479:25]
  wire  arb_io_in_0_ready; // @[Cache.scala 488:19]
  wire  arb_io_in_0_valid; // @[Cache.scala 488:19]
  wire [31:0] arb_io_in_0_bits_addr; // @[Cache.scala 488:19]
  wire [2:0] arb_io_in_0_bits_size; // @[Cache.scala 488:19]
  wire [3:0] arb_io_in_0_bits_cmd; // @[Cache.scala 488:19]
  wire [7:0] arb_io_in_0_bits_wmask; // @[Cache.scala 488:19]
  wire [63:0] arb_io_in_0_bits_wdata; // @[Cache.scala 488:19]
  wire  arb_io_in_1_ready; // @[Cache.scala 488:19]
  wire  arb_io_in_1_valid; // @[Cache.scala 488:19]
  wire [31:0] arb_io_in_1_bits_addr; // @[Cache.scala 488:19]
  wire [2:0] arb_io_in_1_bits_size; // @[Cache.scala 488:19]
  wire [3:0] arb_io_in_1_bits_cmd; // @[Cache.scala 488:19]
  wire [7:0] arb_io_in_1_bits_wmask; // @[Cache.scala 488:19]
  wire [63:0] arb_io_in_1_bits_wdata; // @[Cache.scala 488:19]
  wire  arb_io_out_ready; // @[Cache.scala 488:19]
  wire  arb_io_out_valid; // @[Cache.scala 488:19]
  wire [31:0] arb_io_out_bits_addr; // @[Cache.scala 488:19]
  wire [2:0] arb_io_out_bits_size; // @[Cache.scala 488:19]
  wire [3:0] arb_io_out_bits_cmd; // @[Cache.scala 488:19]
  wire [7:0] arb_io_out_bits_wmask; // @[Cache.scala 488:19]
  wire [63:0] arb_io_out_bits_wdata; // @[Cache.scala 488:19]
  wire  _T = s2_io_out_ready & s2_io_out_valid; // @[Decoupled.scala 40:37]
  reg  _T_2; // @[Pipeline.scala 24:24]
  wire  _GEN_0 = _T ? 1'h0 : _T_2; // @[Pipeline.scala 25:25]
  wire  _T_3 = s1_io_out_valid & s2_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_1 = _T_3 | _GEN_0; // @[Pipeline.scala 26:38]
  reg [31:0] _T_5_req_addr; // @[Reg.scala 15:16]
  reg [2:0] _T_5_req_size; // @[Reg.scala 15:16]
  reg [3:0] _T_5_req_cmd; // @[Reg.scala 15:16]
  reg [7:0] _T_5_req_wmask; // @[Reg.scala 15:16]
  reg [63:0] _T_5_req_wdata; // @[Reg.scala 15:16]
  reg  _T_7; // @[Pipeline.scala 24:24]
  wire  _GEN_8 = s3_io_isFinish ? 1'h0 : _T_7; // @[Pipeline.scala 25:25]
  wire  _T_8 = s2_io_out_valid & s3_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_9 = _T_8 | _GEN_8; // @[Pipeline.scala 26:38]
  reg [31:0] _T_10_req_addr; // @[Reg.scala 15:16]
  reg [2:0] _T_10_req_size; // @[Reg.scala 15:16]
  reg [3:0] _T_10_req_cmd; // @[Reg.scala 15:16]
  reg [7:0] _T_10_req_wmask; // @[Reg.scala 15:16]
  reg [63:0] _T_10_req_wdata; // @[Reg.scala 15:16]
  reg [18:0] _T_10_metas_0_tag; // @[Reg.scala 15:16]
  reg  _T_10_metas_0_valid; // @[Reg.scala 15:16]
  reg  _T_10_metas_0_dirty; // @[Reg.scala 15:16]
  reg [18:0] _T_10_metas_1_tag; // @[Reg.scala 15:16]
  reg  _T_10_metas_1_valid; // @[Reg.scala 15:16]
  reg  _T_10_metas_1_dirty; // @[Reg.scala 15:16]
  reg [18:0] _T_10_metas_2_tag; // @[Reg.scala 15:16]
  reg  _T_10_metas_2_valid; // @[Reg.scala 15:16]
  reg  _T_10_metas_2_dirty; // @[Reg.scala 15:16]
  reg [18:0] _T_10_metas_3_tag; // @[Reg.scala 15:16]
  reg  _T_10_metas_3_valid; // @[Reg.scala 15:16]
  reg  _T_10_metas_3_dirty; // @[Reg.scala 15:16]
  reg [63:0] _T_10_datas_0_data; // @[Reg.scala 15:16]
  reg [63:0] _T_10_datas_1_data; // @[Reg.scala 15:16]
  reg [63:0] _T_10_datas_2_data; // @[Reg.scala 15:16]
  reg [63:0] _T_10_datas_3_data; // @[Reg.scala 15:16]
  reg  _T_10_hit; // @[Reg.scala 15:16]
  reg [3:0] _T_10_waymask; // @[Reg.scala 15:16]
  reg  _T_10_mmio; // @[Reg.scala 15:16]
  reg  _T_10_isForwardData; // @[Reg.scala 15:16]
  reg [63:0] _T_10_forwardData_data_data; // @[Reg.scala 15:16]
  reg [3:0] _T_10_forwardData_waymask; // @[Reg.scala 15:16]
  wire  _T_12 = ~s2_io_in_valid; // @[Cache.scala 503:15]
  wire  _T_13 = ~s3_io_in_valid; // @[Cache.scala 503:34]
  wire  _T_15 = s3_io_out_bits_cmd == 4'h4; // @[SimpleBus.scala 95:26]
  wire  _T_16 = s3_io_out_valid & _T_15; // @[Cache.scala 505:43]
  wire  _T_17 = s3_io_out_valid | s3_io_dataReadRespToL1; // @[Cache.scala 505:100]
  reg [63:0] _T_20; // @[GTimer.scala 24:20]
  wire [63:0] _T_22 = _T_20 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_26 = ~reset; // @[Debug.scala 56:24]
  reg [63:0] _T_29; // @[GTimer.scala 24:20]
  wire [63:0] _T_31 = _T_29 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_38; // @[GTimer.scala 24:20]
  wire [63:0] _T_40 = _T_38 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_47; // @[GTimer.scala 24:20]
  wire [63:0] _T_49 = _T_47 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_56; // @[GTimer.scala 24:20]
  wire [63:0] _T_58 = _T_56 + 64'h1; // @[GTimer.scala 25:12]
  wire  _GEN_39 = s1_io_in_valid & DISPLAY_ENABLE; // @[Debug.scala 56:24]
  wire  _GEN_41 = s2_io_in_valid & DISPLAY_ENABLE; // @[Debug.scala 56:24]
  wire  _GEN_43 = s3_io_in_valid & DISPLAY_ENABLE; // @[Debug.scala 56:24]
  CacheStage1_1 s1 ( // @[Cache.scala 475:18]
    .clock(s1_clock),
    .reset(s1_reset),
    .io_in_ready(s1_io_in_ready),
    .io_in_valid(s1_io_in_valid),
    .io_in_bits_addr(s1_io_in_bits_addr),
    .io_in_bits_size(s1_io_in_bits_size),
    .io_in_bits_cmd(s1_io_in_bits_cmd),
    .io_in_bits_wmask(s1_io_in_bits_wmask),
    .io_in_bits_wdata(s1_io_in_bits_wdata),
    .io_out_ready(s1_io_out_ready),
    .io_out_valid(s1_io_out_valid),
    .io_out_bits_req_addr(s1_io_out_bits_req_addr),
    .io_out_bits_req_size(s1_io_out_bits_req_size),
    .io_out_bits_req_cmd(s1_io_out_bits_req_cmd),
    .io_out_bits_req_wmask(s1_io_out_bits_req_wmask),
    .io_out_bits_req_wdata(s1_io_out_bits_req_wdata),
    .io_metaReadBus_req_ready(s1_io_metaReadBus_req_ready),
    .io_metaReadBus_req_valid(s1_io_metaReadBus_req_valid),
    .io_metaReadBus_req_bits_setIdx(s1_io_metaReadBus_req_bits_setIdx),
    .io_metaReadBus_resp_data_0_tag(s1_io_metaReadBus_resp_data_0_tag),
    .io_metaReadBus_resp_data_0_valid(s1_io_metaReadBus_resp_data_0_valid),
    .io_metaReadBus_resp_data_0_dirty(s1_io_metaReadBus_resp_data_0_dirty),
    .io_metaReadBus_resp_data_1_tag(s1_io_metaReadBus_resp_data_1_tag),
    .io_metaReadBus_resp_data_1_valid(s1_io_metaReadBus_resp_data_1_valid),
    .io_metaReadBus_resp_data_1_dirty(s1_io_metaReadBus_resp_data_1_dirty),
    .io_metaReadBus_resp_data_2_tag(s1_io_metaReadBus_resp_data_2_tag),
    .io_metaReadBus_resp_data_2_valid(s1_io_metaReadBus_resp_data_2_valid),
    .io_metaReadBus_resp_data_2_dirty(s1_io_metaReadBus_resp_data_2_dirty),
    .io_metaReadBus_resp_data_3_tag(s1_io_metaReadBus_resp_data_3_tag),
    .io_metaReadBus_resp_data_3_valid(s1_io_metaReadBus_resp_data_3_valid),
    .io_metaReadBus_resp_data_3_dirty(s1_io_metaReadBus_resp_data_3_dirty),
    .io_dataReadBus_req_ready(s1_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s1_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s1_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s1_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s1_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s1_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s1_io_dataReadBus_resp_data_3_data),
    .DISPLAY_ENABLE(s1_DISPLAY_ENABLE)
  );
  CacheStage2_1 s2 ( // @[Cache.scala 476:18]
    .clock(s2_clock),
    .reset(s2_reset),
    .io_in_ready(s2_io_in_ready),
    .io_in_valid(s2_io_in_valid),
    .io_in_bits_req_addr(s2_io_in_bits_req_addr),
    .io_in_bits_req_size(s2_io_in_bits_req_size),
    .io_in_bits_req_cmd(s2_io_in_bits_req_cmd),
    .io_in_bits_req_wmask(s2_io_in_bits_req_wmask),
    .io_in_bits_req_wdata(s2_io_in_bits_req_wdata),
    .io_out_ready(s2_io_out_ready),
    .io_out_valid(s2_io_out_valid),
    .io_out_bits_req_addr(s2_io_out_bits_req_addr),
    .io_out_bits_req_size(s2_io_out_bits_req_size),
    .io_out_bits_req_cmd(s2_io_out_bits_req_cmd),
    .io_out_bits_req_wmask(s2_io_out_bits_req_wmask),
    .io_out_bits_req_wdata(s2_io_out_bits_req_wdata),
    .io_out_bits_metas_0_tag(s2_io_out_bits_metas_0_tag),
    .io_out_bits_metas_0_valid(s2_io_out_bits_metas_0_valid),
    .io_out_bits_metas_0_dirty(s2_io_out_bits_metas_0_dirty),
    .io_out_bits_metas_1_tag(s2_io_out_bits_metas_1_tag),
    .io_out_bits_metas_1_valid(s2_io_out_bits_metas_1_valid),
    .io_out_bits_metas_1_dirty(s2_io_out_bits_metas_1_dirty),
    .io_out_bits_metas_2_tag(s2_io_out_bits_metas_2_tag),
    .io_out_bits_metas_2_valid(s2_io_out_bits_metas_2_valid),
    .io_out_bits_metas_2_dirty(s2_io_out_bits_metas_2_dirty),
    .io_out_bits_metas_3_tag(s2_io_out_bits_metas_3_tag),
    .io_out_bits_metas_3_valid(s2_io_out_bits_metas_3_valid),
    .io_out_bits_metas_3_dirty(s2_io_out_bits_metas_3_dirty),
    .io_out_bits_datas_0_data(s2_io_out_bits_datas_0_data),
    .io_out_bits_datas_1_data(s2_io_out_bits_datas_1_data),
    .io_out_bits_datas_2_data(s2_io_out_bits_datas_2_data),
    .io_out_bits_datas_3_data(s2_io_out_bits_datas_3_data),
    .io_out_bits_hit(s2_io_out_bits_hit),
    .io_out_bits_waymask(s2_io_out_bits_waymask),
    .io_out_bits_mmio(s2_io_out_bits_mmio),
    .io_out_bits_isForwardData(s2_io_out_bits_isForwardData),
    .io_out_bits_forwardData_data_data(s2_io_out_bits_forwardData_data_data),
    .io_out_bits_forwardData_waymask(s2_io_out_bits_forwardData_waymask),
    .io_metaReadResp_0_tag(s2_io_metaReadResp_0_tag),
    .io_metaReadResp_0_valid(s2_io_metaReadResp_0_valid),
    .io_metaReadResp_0_dirty(s2_io_metaReadResp_0_dirty),
    .io_metaReadResp_1_tag(s2_io_metaReadResp_1_tag),
    .io_metaReadResp_1_valid(s2_io_metaReadResp_1_valid),
    .io_metaReadResp_1_dirty(s2_io_metaReadResp_1_dirty),
    .io_metaReadResp_2_tag(s2_io_metaReadResp_2_tag),
    .io_metaReadResp_2_valid(s2_io_metaReadResp_2_valid),
    .io_metaReadResp_2_dirty(s2_io_metaReadResp_2_dirty),
    .io_metaReadResp_3_tag(s2_io_metaReadResp_3_tag),
    .io_metaReadResp_3_valid(s2_io_metaReadResp_3_valid),
    .io_metaReadResp_3_dirty(s2_io_metaReadResp_3_dirty),
    .io_dataReadResp_0_data(s2_io_dataReadResp_0_data),
    .io_dataReadResp_1_data(s2_io_dataReadResp_1_data),
    .io_dataReadResp_2_data(s2_io_dataReadResp_2_data),
    .io_dataReadResp_3_data(s2_io_dataReadResp_3_data),
    .io_metaWriteBus_req_valid(s2_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s2_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s2_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_data_dirty(s2_io_metaWriteBus_req_bits_data_dirty),
    .io_metaWriteBus_req_bits_waymask(s2_io_metaWriteBus_req_bits_waymask),
    .io_dataWriteBus_req_valid(s2_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s2_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s2_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s2_io_dataWriteBus_req_bits_waymask),
    .DISPLAY_ENABLE(s2_DISPLAY_ENABLE)
  );
  CacheStage3_1 s3 ( // @[Cache.scala 477:18]
    .clock(s3_clock),
    .reset(s3_reset),
    .io_in_ready(s3_io_in_ready),
    .io_in_valid(s3_io_in_valid),
    .io_in_bits_req_addr(s3_io_in_bits_req_addr),
    .io_in_bits_req_size(s3_io_in_bits_req_size),
    .io_in_bits_req_cmd(s3_io_in_bits_req_cmd),
    .io_in_bits_req_wmask(s3_io_in_bits_req_wmask),
    .io_in_bits_req_wdata(s3_io_in_bits_req_wdata),
    .io_in_bits_metas_0_tag(s3_io_in_bits_metas_0_tag),
    .io_in_bits_metas_0_valid(s3_io_in_bits_metas_0_valid),
    .io_in_bits_metas_0_dirty(s3_io_in_bits_metas_0_dirty),
    .io_in_bits_metas_1_tag(s3_io_in_bits_metas_1_tag),
    .io_in_bits_metas_1_valid(s3_io_in_bits_metas_1_valid),
    .io_in_bits_metas_1_dirty(s3_io_in_bits_metas_1_dirty),
    .io_in_bits_metas_2_tag(s3_io_in_bits_metas_2_tag),
    .io_in_bits_metas_2_valid(s3_io_in_bits_metas_2_valid),
    .io_in_bits_metas_2_dirty(s3_io_in_bits_metas_2_dirty),
    .io_in_bits_metas_3_tag(s3_io_in_bits_metas_3_tag),
    .io_in_bits_metas_3_valid(s3_io_in_bits_metas_3_valid),
    .io_in_bits_metas_3_dirty(s3_io_in_bits_metas_3_dirty),
    .io_in_bits_datas_0_data(s3_io_in_bits_datas_0_data),
    .io_in_bits_datas_1_data(s3_io_in_bits_datas_1_data),
    .io_in_bits_datas_2_data(s3_io_in_bits_datas_2_data),
    .io_in_bits_datas_3_data(s3_io_in_bits_datas_3_data),
    .io_in_bits_hit(s3_io_in_bits_hit),
    .io_in_bits_waymask(s3_io_in_bits_waymask),
    .io_in_bits_mmio(s3_io_in_bits_mmio),
    .io_in_bits_isForwardData(s3_io_in_bits_isForwardData),
    .io_in_bits_forwardData_data_data(s3_io_in_bits_forwardData_data_data),
    .io_in_bits_forwardData_waymask(s3_io_in_bits_forwardData_waymask),
    .io_out_ready(s3_io_out_ready),
    .io_out_valid(s3_io_out_valid),
    .io_out_bits_cmd(s3_io_out_bits_cmd),
    .io_out_bits_rdata(s3_io_out_bits_rdata),
    .io_isFinish(s3_io_isFinish),
    .io_dataReadBus_req_ready(s3_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s3_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s3_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s3_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s3_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s3_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s3_io_dataReadBus_resp_data_3_data),
    .io_dataWriteBus_req_valid(s3_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s3_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s3_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s3_io_dataWriteBus_req_bits_waymask),
    .io_metaWriteBus_req_valid(s3_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s3_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s3_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_data_valid(s3_io_metaWriteBus_req_bits_data_valid),
    .io_metaWriteBus_req_bits_data_dirty(s3_io_metaWriteBus_req_bits_data_dirty),
    .io_metaWriteBus_req_bits_waymask(s3_io_metaWriteBus_req_bits_waymask),
    .io_mem_req_ready(s3_io_mem_req_ready),
    .io_mem_req_valid(s3_io_mem_req_valid),
    .io_mem_req_bits_addr(s3_io_mem_req_bits_addr),
    .io_mem_req_bits_size(s3_io_mem_req_bits_size),
    .io_mem_req_bits_cmd(s3_io_mem_req_bits_cmd),
    .io_mem_req_bits_wmask(s3_io_mem_req_bits_wmask),
    .io_mem_req_bits_wdata(s3_io_mem_req_bits_wdata),
    .io_mem_resp_ready(s3_io_mem_resp_ready),
    .io_mem_resp_valid(s3_io_mem_resp_valid),
    .io_mem_resp_bits_cmd(s3_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_rdata(s3_io_mem_resp_bits_rdata),
    .io_mmio_req_ready(s3_io_mmio_req_ready),
    .io_mmio_req_valid(s3_io_mmio_req_valid),
    .io_mmio_req_bits_addr(s3_io_mmio_req_bits_addr),
    .io_mmio_req_bits_size(s3_io_mmio_req_bits_size),
    .io_mmio_req_bits_cmd(s3_io_mmio_req_bits_cmd),
    .io_mmio_req_bits_wmask(s3_io_mmio_req_bits_wmask),
    .io_mmio_req_bits_wdata(s3_io_mmio_req_bits_wdata),
    .io_mmio_resp_ready(s3_io_mmio_resp_ready),
    .io_mmio_resp_valid(s3_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(s3_io_mmio_resp_bits_rdata),
    .io_cohResp_valid(s3_io_cohResp_valid),
    .io_cohResp_bits_cmd(s3_io_cohResp_bits_cmd),
    .io_cohResp_bits_rdata(s3_io_cohResp_bits_rdata),
    .io_dataReadRespToL1(s3_io_dataReadRespToL1),
    .mmio_0(s3_mmio_0),
    .DISPLAY_ENABLE(s3_DISPLAY_ENABLE)
  );
  SRAMTemplateWithArbiter metaArray ( // @[Cache.scala 478:25]
    .clock(metaArray_clock),
    .reset(metaArray_reset),
    .io_r_0_req_ready(metaArray_io_r_0_req_ready),
    .io_r_0_req_valid(metaArray_io_r_0_req_valid),
    .io_r_0_req_bits_setIdx(metaArray_io_r_0_req_bits_setIdx),
    .io_r_0_resp_data_0_tag(metaArray_io_r_0_resp_data_0_tag),
    .io_r_0_resp_data_0_valid(metaArray_io_r_0_resp_data_0_valid),
    .io_r_0_resp_data_0_dirty(metaArray_io_r_0_resp_data_0_dirty),
    .io_r_0_resp_data_1_tag(metaArray_io_r_0_resp_data_1_tag),
    .io_r_0_resp_data_1_valid(metaArray_io_r_0_resp_data_1_valid),
    .io_r_0_resp_data_1_dirty(metaArray_io_r_0_resp_data_1_dirty),
    .io_r_0_resp_data_2_tag(metaArray_io_r_0_resp_data_2_tag),
    .io_r_0_resp_data_2_valid(metaArray_io_r_0_resp_data_2_valid),
    .io_r_0_resp_data_2_dirty(metaArray_io_r_0_resp_data_2_dirty),
    .io_r_0_resp_data_3_tag(metaArray_io_r_0_resp_data_3_tag),
    .io_r_0_resp_data_3_valid(metaArray_io_r_0_resp_data_3_valid),
    .io_r_0_resp_data_3_dirty(metaArray_io_r_0_resp_data_3_dirty),
    .io_w_req_valid(metaArray_io_w_req_valid),
    .io_w_req_bits_setIdx(metaArray_io_w_req_bits_setIdx),
    .io_w_req_bits_data_tag(metaArray_io_w_req_bits_data_tag),
    .io_w_req_bits_data_dirty(metaArray_io_w_req_bits_data_dirty),
    .io_w_req_bits_waymask(metaArray_io_w_req_bits_waymask)
  );
  SRAMTemplateWithArbiter_1 dataArray ( // @[Cache.scala 479:25]
    .clock(dataArray_clock),
    .reset(dataArray_reset),
    .io_r_0_req_ready(dataArray_io_r_0_req_ready),
    .io_r_0_req_valid(dataArray_io_r_0_req_valid),
    .io_r_0_req_bits_setIdx(dataArray_io_r_0_req_bits_setIdx),
    .io_r_0_resp_data_0_data(dataArray_io_r_0_resp_data_0_data),
    .io_r_0_resp_data_1_data(dataArray_io_r_0_resp_data_1_data),
    .io_r_0_resp_data_2_data(dataArray_io_r_0_resp_data_2_data),
    .io_r_0_resp_data_3_data(dataArray_io_r_0_resp_data_3_data),
    .io_r_1_req_ready(dataArray_io_r_1_req_ready),
    .io_r_1_req_valid(dataArray_io_r_1_req_valid),
    .io_r_1_req_bits_setIdx(dataArray_io_r_1_req_bits_setIdx),
    .io_r_1_resp_data_0_data(dataArray_io_r_1_resp_data_0_data),
    .io_r_1_resp_data_1_data(dataArray_io_r_1_resp_data_1_data),
    .io_r_1_resp_data_2_data(dataArray_io_r_1_resp_data_2_data),
    .io_r_1_resp_data_3_data(dataArray_io_r_1_resp_data_3_data),
    .io_w_req_valid(dataArray_io_w_req_valid),
    .io_w_req_bits_setIdx(dataArray_io_w_req_bits_setIdx),
    .io_w_req_bits_data_data(dataArray_io_w_req_bits_data_data),
    .io_w_req_bits_waymask(dataArray_io_w_req_bits_waymask)
  );
  Arbiter_9 arb ( // @[Cache.scala 488:19]
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_addr(arb_io_in_0_bits_addr),
    .io_in_0_bits_size(arb_io_in_0_bits_size),
    .io_in_0_bits_cmd(arb_io_in_0_bits_cmd),
    .io_in_0_bits_wmask(arb_io_in_0_bits_wmask),
    .io_in_0_bits_wdata(arb_io_in_0_bits_wdata),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_addr(arb_io_in_1_bits_addr),
    .io_in_1_bits_size(arb_io_in_1_bits_size),
    .io_in_1_bits_cmd(arb_io_in_1_bits_cmd),
    .io_in_1_bits_wmask(arb_io_in_1_bits_wmask),
    .io_in_1_bits_wdata(arb_io_in_1_bits_wdata),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_addr(arb_io_out_bits_addr),
    .io_out_bits_size(arb_io_out_bits_size),
    .io_out_bits_cmd(arb_io_out_bits_cmd),
    .io_out_bits_wmask(arb_io_out_bits_wmask),
    .io_out_bits_wdata(arb_io_out_bits_wdata)
  );
  assign io_in_req_ready = arb_io_in_1_ready; // @[Cache.scala 489:28]
  assign io_in_resp_valid = _T_16 ? 1'h0 : _T_17; // @[Cache.scala 499:14 Cache.scala 505:20]
  assign io_in_resp_bits_cmd = s3_io_out_bits_cmd; // @[Cache.scala 499:14]
  assign io_in_resp_bits_rdata = s3_io_out_bits_rdata; // @[Cache.scala 499:14]
  assign io_out_mem_req_valid = s3_io_mem_req_valid; // @[Cache.scala 501:14]
  assign io_out_mem_req_bits_addr = s3_io_mem_req_bits_addr; // @[Cache.scala 501:14]
  assign io_out_mem_req_bits_cmd = s3_io_mem_req_bits_cmd; // @[Cache.scala 501:14]
  assign io_out_mem_req_bits_wdata = s3_io_mem_req_bits_wdata; // @[Cache.scala 501:14]
  assign io_out_coh_req_ready = arb_io_in_0_ready; // @[Cache.scala 514:26]
  assign io_out_coh_resp_valid = s3_io_cohResp_valid; // @[Cache.scala 515:21]
  assign io_out_coh_resp_bits_cmd = s3_io_cohResp_bits_cmd; // @[Cache.scala 515:21]
  assign io_out_coh_resp_bits_rdata = s3_io_cohResp_bits_rdata; // @[Cache.scala 515:21]
  assign io_mmio_req_valid = s3_io_mmio_req_valid; // @[Cache.scala 502:11]
  assign io_mmio_req_bits_addr = s3_io_mmio_req_bits_addr; // @[Cache.scala 502:11]
  assign io_mmio_req_bits_size = s3_io_mmio_req_bits_size; // @[Cache.scala 502:11]
  assign io_mmio_req_bits_cmd = s3_io_mmio_req_bits_cmd; // @[Cache.scala 502:11]
  assign io_mmio_req_bits_wmask = s3_io_mmio_req_bits_wmask; // @[Cache.scala 502:11]
  assign io_mmio_req_bits_wdata = s3_io_mmio_req_bits_wdata; // @[Cache.scala 502:11]
  assign io_empty = _T_12 & _T_13; // @[Cache.scala 503:12]
  assign mmio = s3_mmio_0;
  assign s1_clock = clock;
  assign s1_reset = reset;
  assign s1_io_in_valid = arb_io_out_valid; // @[Cache.scala 491:12]
  assign s1_io_in_bits_addr = arb_io_out_bits_addr; // @[Cache.scala 491:12]
  assign s1_io_in_bits_size = arb_io_out_bits_size; // @[Cache.scala 491:12]
  assign s1_io_in_bits_cmd = arb_io_out_bits_cmd; // @[Cache.scala 491:12]
  assign s1_io_in_bits_wmask = arb_io_out_bits_wmask; // @[Cache.scala 491:12]
  assign s1_io_in_bits_wdata = arb_io_out_bits_wdata; // @[Cache.scala 491:12]
  assign s1_io_out_ready = s2_io_in_ready; // @[Pipeline.scala 29:16]
  assign s1_io_metaReadBus_req_ready = metaArray_io_r_0_req_ready; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_0_tag = metaArray_io_r_0_resp_data_0_tag; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_0_valid = metaArray_io_r_0_resp_data_0_valid; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_0_dirty = metaArray_io_r_0_resp_data_0_dirty; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_1_tag = metaArray_io_r_0_resp_data_1_tag; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_1_valid = metaArray_io_r_0_resp_data_1_valid; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_1_dirty = metaArray_io_r_0_resp_data_1_dirty; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_2_tag = metaArray_io_r_0_resp_data_2_tag; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_2_valid = metaArray_io_r_0_resp_data_2_valid; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_2_dirty = metaArray_io_r_0_resp_data_2_dirty; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_3_tag = metaArray_io_r_0_resp_data_3_tag; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_3_valid = metaArray_io_r_0_resp_data_3_valid; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_3_dirty = metaArray_io_r_0_resp_data_3_dirty; // @[Cache.scala 523:21]
  assign s1_io_dataReadBus_req_ready = dataArray_io_r_0_req_ready; // @[Cache.scala 524:21]
  assign s1_io_dataReadBus_resp_data_0_data = dataArray_io_r_0_resp_data_0_data; // @[Cache.scala 524:21]
  assign s1_io_dataReadBus_resp_data_1_data = dataArray_io_r_0_resp_data_1_data; // @[Cache.scala 524:21]
  assign s1_io_dataReadBus_resp_data_2_data = dataArray_io_r_0_resp_data_2_data; // @[Cache.scala 524:21]
  assign s1_io_dataReadBus_resp_data_3_data = dataArray_io_r_0_resp_data_3_data; // @[Cache.scala 524:21]
  assign s1_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign s2_clock = clock;
  assign s2_reset = reset;
  assign s2_io_in_valid = _T_2; // @[Pipeline.scala 31:17]
  assign s2_io_in_bits_req_addr = _T_5_req_addr; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_size = _T_5_req_size; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_cmd = _T_5_req_cmd; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_wmask = _T_5_req_wmask; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_wdata = _T_5_req_wdata; // @[Pipeline.scala 30:16]
  assign s2_io_out_ready = s3_io_in_ready; // @[Pipeline.scala 29:16]
  assign s2_io_metaReadResp_0_tag = s1_io_metaReadBus_resp_data_0_tag; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_0_valid = s1_io_metaReadBus_resp_data_0_valid; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_0_dirty = s1_io_metaReadBus_resp_data_0_dirty; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_1_tag = s1_io_metaReadBus_resp_data_1_tag; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_1_valid = s1_io_metaReadBus_resp_data_1_valid; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_1_dirty = s1_io_metaReadBus_resp_data_1_dirty; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_2_tag = s1_io_metaReadBus_resp_data_2_tag; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_2_valid = s1_io_metaReadBus_resp_data_2_valid; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_2_dirty = s1_io_metaReadBus_resp_data_2_dirty; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_3_tag = s1_io_metaReadBus_resp_data_3_tag; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_3_valid = s1_io_metaReadBus_resp_data_3_valid; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_3_dirty = s1_io_metaReadBus_resp_data_3_dirty; // @[Cache.scala 530:22]
  assign s2_io_dataReadResp_0_data = s1_io_dataReadBus_resp_data_0_data; // @[Cache.scala 531:22]
  assign s2_io_dataReadResp_1_data = s1_io_dataReadBus_resp_data_1_data; // @[Cache.scala 531:22]
  assign s2_io_dataReadResp_2_data = s1_io_dataReadBus_resp_data_2_data; // @[Cache.scala 531:22]
  assign s2_io_dataReadResp_3_data = s1_io_dataReadBus_resp_data_3_data; // @[Cache.scala 531:22]
  assign s2_io_metaWriteBus_req_valid = s3_io_metaWriteBus_req_valid; // @[Cache.scala 533:22]
  assign s2_io_metaWriteBus_req_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 533:22]
  assign s2_io_metaWriteBus_req_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 533:22]
  assign s2_io_metaWriteBus_req_bits_data_dirty = s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 533:22]
  assign s2_io_metaWriteBus_req_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 533:22]
  assign s2_io_dataWriteBus_req_valid = s3_io_dataWriteBus_req_valid; // @[Cache.scala 532:22]
  assign s2_io_dataWriteBus_req_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 532:22]
  assign s2_io_dataWriteBus_req_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 532:22]
  assign s2_io_dataWriteBus_req_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 532:22]
  assign s2_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign s3_clock = clock;
  assign s3_reset = reset;
  assign s3_io_in_valid = _T_7; // @[Pipeline.scala 31:17]
  assign s3_io_in_bits_req_addr = _T_10_req_addr; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_size = _T_10_req_size; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_cmd = _T_10_req_cmd; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_wmask = _T_10_req_wmask; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_wdata = _T_10_req_wdata; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_tag = _T_10_metas_0_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_valid = _T_10_metas_0_valid; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_dirty = _T_10_metas_0_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_tag = _T_10_metas_1_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_valid = _T_10_metas_1_valid; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_dirty = _T_10_metas_1_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_tag = _T_10_metas_2_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_valid = _T_10_metas_2_valid; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_dirty = _T_10_metas_2_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_tag = _T_10_metas_3_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_valid = _T_10_metas_3_valid; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_dirty = _T_10_metas_3_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_0_data = _T_10_datas_0_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_1_data = _T_10_datas_1_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_2_data = _T_10_datas_2_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_3_data = _T_10_datas_3_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_hit = _T_10_hit; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_waymask = _T_10_waymask; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_mmio = _T_10_mmio; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_isForwardData = _T_10_isForwardData; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_data_data = _T_10_forwardData_data_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_waymask = _T_10_forwardData_waymask; // @[Pipeline.scala 30:16]
  assign s3_io_out_ready = io_in_resp_ready; // @[Cache.scala 499:14]
  assign s3_io_dataReadBus_req_ready = dataArray_io_r_1_req_ready; // @[Cache.scala 525:21]
  assign s3_io_dataReadBus_resp_data_0_data = dataArray_io_r_1_resp_data_0_data; // @[Cache.scala 525:21]
  assign s3_io_dataReadBus_resp_data_1_data = dataArray_io_r_1_resp_data_1_data; // @[Cache.scala 525:21]
  assign s3_io_dataReadBus_resp_data_2_data = dataArray_io_r_1_resp_data_2_data; // @[Cache.scala 525:21]
  assign s3_io_dataReadBus_resp_data_3_data = dataArray_io_r_1_resp_data_3_data; // @[Cache.scala 525:21]
  assign s3_io_mem_req_ready = io_out_mem_req_ready; // @[Cache.scala 501:14]
  assign s3_io_mem_resp_valid = io_out_mem_resp_valid; // @[Cache.scala 501:14]
  assign s3_io_mem_resp_bits_cmd = io_out_mem_resp_bits_cmd; // @[Cache.scala 501:14]
  assign s3_io_mem_resp_bits_rdata = io_out_mem_resp_bits_rdata; // @[Cache.scala 501:14]
  assign s3_io_mmio_req_ready = io_mmio_req_ready; // @[Cache.scala 502:11]
  assign s3_io_mmio_resp_valid = io_mmio_resp_valid; // @[Cache.scala 502:11]
  assign s3_io_mmio_resp_bits_rdata = io_mmio_resp_bits_rdata; // @[Cache.scala 502:11]
  assign s3_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign metaArray_clock = clock;
  assign metaArray_reset = reset;
  assign metaArray_io_r_0_req_valid = s1_io_metaReadBus_req_valid; // @[Cache.scala 523:21]
  assign metaArray_io_r_0_req_bits_setIdx = s1_io_metaReadBus_req_bits_setIdx; // @[Cache.scala 523:21]
  assign metaArray_io_w_req_valid = s3_io_metaWriteBus_req_valid; // @[Cache.scala 527:18]
  assign metaArray_io_w_req_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 527:18]
  assign metaArray_io_w_req_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 527:18]
  assign metaArray_io_w_req_bits_data_dirty = s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 527:18]
  assign metaArray_io_w_req_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 527:18]
  assign dataArray_clock = clock;
  assign dataArray_reset = reset;
  assign dataArray_io_r_0_req_valid = s1_io_dataReadBus_req_valid; // @[Cache.scala 524:21]
  assign dataArray_io_r_0_req_bits_setIdx = s1_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 524:21]
  assign dataArray_io_r_1_req_valid = s3_io_dataReadBus_req_valid; // @[Cache.scala 525:21]
  assign dataArray_io_r_1_req_bits_setIdx = s3_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 525:21]
  assign dataArray_io_w_req_valid = s3_io_dataWriteBus_req_valid; // @[Cache.scala 528:18]
  assign dataArray_io_w_req_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 528:18]
  assign dataArray_io_w_req_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 528:18]
  assign dataArray_io_w_req_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 528:18]
  assign arb_io_in_0_valid = io_out_coh_req_valid; // @[Cache.scala 513:24]
  assign arb_io_in_0_bits_addr = io_out_coh_req_bits_addr; // @[Cache.scala 512:23]
  assign arb_io_in_0_bits_size = 3'h3; // @[Cache.scala 512:23]
  assign arb_io_in_0_bits_cmd = 4'h8; // @[Cache.scala 512:23]
  assign arb_io_in_0_bits_wmask = 8'hff; // @[Cache.scala 512:23]
  assign arb_io_in_0_bits_wdata = io_out_coh_req_bits_wdata; // @[Cache.scala 512:23]
  assign arb_io_in_1_valid = io_in_req_valid; // @[Cache.scala 489:28]
  assign arb_io_in_1_bits_addr = io_in_req_bits_addr; // @[Cache.scala 489:28]
  assign arb_io_in_1_bits_size = io_in_req_bits_size; // @[Cache.scala 489:28]
  assign arb_io_in_1_bits_cmd = io_in_req_bits_cmd; // @[Cache.scala 489:28]
  assign arb_io_in_1_bits_wmask = io_in_req_bits_wmask; // @[Cache.scala 489:28]
  assign arb_io_in_1_bits_wdata = io_in_req_bits_wdata; // @[Cache.scala 489:28]
  assign arb_io_out_ready = s1_io_in_ready; // @[Cache.scala 491:12]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _T_5_req_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_5_req_size = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  _T_5_req_cmd = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  _T_5_req_wmask = _RAND_4[7:0];
  _RAND_5 = {2{`RANDOM}};
  _T_5_req_wdata = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  _T_7 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_10_req_addr = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  _T_10_req_size = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  _T_10_req_cmd = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  _T_10_req_wmask = _RAND_10[7:0];
  _RAND_11 = {2{`RANDOM}};
  _T_10_req_wdata = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  _T_10_metas_0_tag = _RAND_12[18:0];
  _RAND_13 = {1{`RANDOM}};
  _T_10_metas_0_valid = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  _T_10_metas_0_dirty = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  _T_10_metas_1_tag = _RAND_15[18:0];
  _RAND_16 = {1{`RANDOM}};
  _T_10_metas_1_valid = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  _T_10_metas_1_dirty = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  _T_10_metas_2_tag = _RAND_18[18:0];
  _RAND_19 = {1{`RANDOM}};
  _T_10_metas_2_valid = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  _T_10_metas_2_dirty = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  _T_10_metas_3_tag = _RAND_21[18:0];
  _RAND_22 = {1{`RANDOM}};
  _T_10_metas_3_valid = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  _T_10_metas_3_dirty = _RAND_23[0:0];
  _RAND_24 = {2{`RANDOM}};
  _T_10_datas_0_data = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  _T_10_datas_1_data = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  _T_10_datas_2_data = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  _T_10_datas_3_data = _RAND_27[63:0];
  _RAND_28 = {1{`RANDOM}};
  _T_10_hit = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  _T_10_waymask = _RAND_29[3:0];
  _RAND_30 = {1{`RANDOM}};
  _T_10_mmio = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  _T_10_isForwardData = _RAND_31[0:0];
  _RAND_32 = {2{`RANDOM}};
  _T_10_forwardData_data_data = _RAND_32[63:0];
  _RAND_33 = {1{`RANDOM}};
  _T_10_forwardData_waymask = _RAND_33[3:0];
  _RAND_34 = {2{`RANDOM}};
  _T_20 = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  _T_29 = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  _T_38 = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  _T_47 = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  _T_56 = _RAND_38[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_2 <= 1'h0;
    end else begin
      _T_2 <= _GEN_1;
    end
    if (_T_3) begin
      _T_5_req_addr <= s1_io_out_bits_req_addr;
    end
    if (_T_3) begin
      _T_5_req_size <= s1_io_out_bits_req_size;
    end
    if (_T_3) begin
      _T_5_req_cmd <= s1_io_out_bits_req_cmd;
    end
    if (_T_3) begin
      _T_5_req_wmask <= s1_io_out_bits_req_wmask;
    end
    if (_T_3) begin
      _T_5_req_wdata <= s1_io_out_bits_req_wdata;
    end
    if (reset) begin
      _T_7 <= 1'h0;
    end else begin
      _T_7 <= _GEN_9;
    end
    if (_T_8) begin
      _T_10_req_addr <= s2_io_out_bits_req_addr;
    end
    if (_T_8) begin
      _T_10_req_size <= s2_io_out_bits_req_size;
    end
    if (_T_8) begin
      _T_10_req_cmd <= s2_io_out_bits_req_cmd;
    end
    if (_T_8) begin
      _T_10_req_wmask <= s2_io_out_bits_req_wmask;
    end
    if (_T_8) begin
      _T_10_req_wdata <= s2_io_out_bits_req_wdata;
    end
    if (_T_8) begin
      _T_10_metas_0_tag <= s2_io_out_bits_metas_0_tag;
    end
    if (_T_8) begin
      _T_10_metas_0_valid <= s2_io_out_bits_metas_0_valid;
    end
    if (_T_8) begin
      _T_10_metas_0_dirty <= s2_io_out_bits_metas_0_dirty;
    end
    if (_T_8) begin
      _T_10_metas_1_tag <= s2_io_out_bits_metas_1_tag;
    end
    if (_T_8) begin
      _T_10_metas_1_valid <= s2_io_out_bits_metas_1_valid;
    end
    if (_T_8) begin
      _T_10_metas_1_dirty <= s2_io_out_bits_metas_1_dirty;
    end
    if (_T_8) begin
      _T_10_metas_2_tag <= s2_io_out_bits_metas_2_tag;
    end
    if (_T_8) begin
      _T_10_metas_2_valid <= s2_io_out_bits_metas_2_valid;
    end
    if (_T_8) begin
      _T_10_metas_2_dirty <= s2_io_out_bits_metas_2_dirty;
    end
    if (_T_8) begin
      _T_10_metas_3_tag <= s2_io_out_bits_metas_3_tag;
    end
    if (_T_8) begin
      _T_10_metas_3_valid <= s2_io_out_bits_metas_3_valid;
    end
    if (_T_8) begin
      _T_10_metas_3_dirty <= s2_io_out_bits_metas_3_dirty;
    end
    if (_T_8) begin
      _T_10_datas_0_data <= s2_io_out_bits_datas_0_data;
    end
    if (_T_8) begin
      _T_10_datas_1_data <= s2_io_out_bits_datas_1_data;
    end
    if (_T_8) begin
      _T_10_datas_2_data <= s2_io_out_bits_datas_2_data;
    end
    if (_T_8) begin
      _T_10_datas_3_data <= s2_io_out_bits_datas_3_data;
    end
    if (_T_8) begin
      _T_10_hit <= s2_io_out_bits_hit;
    end
    if (_T_8) begin
      _T_10_waymask <= s2_io_out_bits_waymask;
    end
    if (_T_8) begin
      _T_10_mmio <= s2_io_out_bits_mmio;
    end
    if (_T_8) begin
      _T_10_isForwardData <= s2_io_out_bits_isForwardData;
    end
    if (_T_8) begin
      _T_10_forwardData_data_data <= s2_io_out_bits_forwardData_data_data;
    end
    if (_T_8) begin
      _T_10_forwardData_waymask <= s2_io_out_bits_forwardData_waymask;
    end
    if (reset) begin
      _T_20 <= 64'h0;
    end else begin
      _T_20 <= _T_22;
    end
    if (reset) begin
      _T_29 <= 64'h0;
    end else begin
      _T_29 <= _T_31;
    end
    if (reset) begin
      _T_38 <= 64'h0;
    end else begin
      _T_38 <= _T_40;
    end
    if (reset) begin
      _T_47 <= 64'h0;
    end else begin
      _T_47 <= _T_49;
    end
    if (reset) begin
      _T_56 <= 64'h0;
    end else begin
      _T_56 <= _T_58;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_26) begin
          $fwrite(32'h80000002,"[%d] Cache_1: ",_T_20); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_26) begin
          $fwrite(32'h80000002,"InReq(%d, %d) InResp(%d, %d) \n",io_in_req_valid,io_in_req_ready,io_in_resp_valid,io_in_resp_ready); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_26) begin
          $fwrite(32'h80000002,"[%d] Cache_1: ",_T_29); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_26) begin
          $fwrite(32'h80000002,"{IN s1:(%d,%d), s2:(%d,%d), s3:(%d,%d)} {OUT s1:(%d,%d), s2:(%d,%d), s3:(%d,%d)}\n",s1_io_in_valid,s1_io_in_ready,s2_io_in_valid,s2_io_in_ready,s3_io_in_valid,s3_io_in_ready,s1_io_out_valid,s1_io_out_ready,s2_io_out_valid,s2_io_out_ready,s3_io_out_valid,s3_io_out_ready); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_39 & _T_26) begin
          $fwrite(32'h80000002,"[%d] Cache_1: ",_T_38); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_39 & _T_26) begin
          $fwrite(32'h80000002,"[dcache.S1]: addr = 0x%x, cmd = %d, size = %d, wmask = 0x%x, wdata = 0x%x\n",s1_io_in_bits_addr,s1_io_in_bits_cmd,s1_io_in_bits_size,s1_io_in_bits_wmask,s1_io_in_bits_wdata); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_26) begin
          $fwrite(32'h80000002,"[%d] Cache_1: ",_T_47); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_26) begin
          $fwrite(32'h80000002,"[dcache.S2]: addr = 0x%x, cmd = %d, size = %d, wmask = 0x%x, wdata = 0x%x\n",s2_io_in_bits_req_addr,s2_io_in_bits_req_cmd,s2_io_in_bits_req_size,s2_io_in_bits_req_wmask,s2_io_in_bits_req_wdata); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_43 & _T_26) begin
          $fwrite(32'h80000002,"[%d] Cache_1: ",_T_56); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_43 & _T_26) begin
          $fwrite(32'h80000002,"[dcache.S3]: addr = 0x%x, cmd = %d, size = %d, wmask = 0x%x, wdata = 0x%x\n",s3_io_in_bits_req_addr,s3_io_in_bits_req_cmd,s3_io_in_bits_req_size,s3_io_in_bits_req_wmask,s3_io_in_bits_req_wdata); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module NutCore(
  input         clock,
  input         reset,
  input         io_imem_mem_req_ready,
  output        io_imem_mem_req_valid,
  output [31:0] io_imem_mem_req_bits_addr,
  output [3:0]  io_imem_mem_req_bits_cmd,
  output [63:0] io_imem_mem_req_bits_wdata,
  input         io_imem_mem_resp_valid,
  input  [3:0]  io_imem_mem_resp_bits_cmd,
  input  [63:0] io_imem_mem_resp_bits_rdata,
  input         io_dmem_mem_req_ready,
  output        io_dmem_mem_req_valid,
  output [31:0] io_dmem_mem_req_bits_addr,
  output [3:0]  io_dmem_mem_req_bits_cmd,
  output [63:0] io_dmem_mem_req_bits_wdata,
  input         io_dmem_mem_resp_valid,
  input  [3:0]  io_dmem_mem_resp_bits_cmd,
  input  [63:0] io_dmem_mem_resp_bits_rdata,
  output        io_dmem_coh_req_ready,
  input         io_dmem_coh_req_valid,
  input  [31:0] io_dmem_coh_req_bits_addr,
  input  [63:0] io_dmem_coh_req_bits_wdata,
  output        io_dmem_coh_resp_valid,
  output [3:0]  io_dmem_coh_resp_bits_cmd,
  output [63:0] io_dmem_coh_resp_bits_rdata,
  input         io_mmio_req_ready,
  output        io_mmio_req_valid,
  output [31:0] io_mmio_req_bits_addr,
  output [2:0]  io_mmio_req_bits_size,
  output [3:0]  io_mmio_req_bits_cmd,
  output [7:0]  io_mmio_req_bits_wmask,
  output [63:0] io_mmio_req_bits_wdata,
  input         io_mmio_resp_valid,
  input  [63:0] io_mmio_resp_bits_rdata,
  output        io_frontend_req_ready,
  input         io_frontend_req_valid,
  input  [31:0] io_frontend_req_bits_addr,
  input  [2:0]  io_frontend_req_bits_size,
  input  [3:0]  io_frontend_req_bits_cmd,
  input  [7:0]  io_frontend_req_bits_wmask,
  input  [63:0] io_frontend_req_bits_wdata,
  input         io_frontend_resp_ready,
  output        io_frontend_resp_valid,
  output [3:0]  io_frontend_resp_bits_cmd,
  output [63:0] io_frontend_resp_bits_rdata,
  output [63:0] _T_4181,
  output [63:0] _T_4184,
  output [63:0] _T_4185,
  output        falseWire,
  output        falseWire_0,
  output [1:0]  _T_4178,
  output [63:0] _T_284_0,
  output [63:0] _T_284_1,
  output [63:0] _T_284_2,
  output [63:0] _T_284_3,
  output [63:0] _T_284_4,
  output [63:0] _T_284_5,
  output [63:0] _T_284_6,
  output [63:0] _T_284_7,
  output [63:0] _T_284_8,
  output [63:0] _T_284_9,
  output [63:0] _T_284_10,
  output [63:0] _T_284_11,
  output [63:0] _T_284_12,
  output [63:0] _T_284_13,
  output [63:0] _T_284_14,
  output [63:0] _T_284_15,
  output [63:0] _T_284_16,
  output [63:0] _T_284_17,
  output [63:0] _T_284_18,
  output [63:0] _T_284_19,
  output [63:0] _T_284_20,
  output [63:0] _T_284_21,
  output [63:0] _T_284_22,
  output [63:0] _T_284_23,
  output [63:0] _T_284_24,
  output [63:0] _T_284_25,
  output [63:0] _T_284_26,
  output [63:0] _T_284_27,
  output [63:0] _T_284_28,
  output [63:0] _T_284_29,
  output [63:0] _T_284_30,
  output [63:0] _T_284_31,
  output        _T_36_0,
  input         io_extra_mtip,
  output [63:0] _T_32_0,
  input         DISPLAY_ENABLE,
  input         io_extra_meip_0,
  output [63:0] _T_31_0,
  output [63:0] _T_37_0,
  output        _T_26_0,
  output        _T_0,
  input         io_extra_msip,
  output [63:0] _T_4183,
  output [63:0] _T_4182,
  output        _T_33_0,
  output [63:0] _T_4179
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [63:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [63:0] _RAND_122;
`endif // RANDOMIZE_REG_INIT
  wire  frontend_clock; // @[NutCore.scala 102:34]
  wire  frontend_reset; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_ready; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_valid; // @[NutCore.scala 102:34]
  wire [63:0] frontend_io_out_0_bits_cf_instr; // @[NutCore.scala 102:34]
  wire [38:0] frontend_io_out_0_bits_cf_pc; // @[NutCore.scala 102:34]
  wire [38:0] frontend_io_out_0_bits_cf_pnpc; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_cf_exceptionVec_1; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_cf_exceptionVec_2; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_cf_exceptionVec_12; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_cf_intrVec_0; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_cf_intrVec_1; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_cf_intrVec_2; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_cf_intrVec_3; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_cf_intrVec_4; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_cf_intrVec_5; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_cf_intrVec_6; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_cf_intrVec_7; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_cf_intrVec_8; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_cf_intrVec_9; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_cf_intrVec_10; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_cf_intrVec_11; // @[NutCore.scala 102:34]
  wire [3:0] frontend_io_out_0_bits_cf_brIdx; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_cf_crossPageIPFFix; // @[NutCore.scala 102:34]
  wire [1:0] frontend_io_out_0_bits_ctrl_src1Type; // @[NutCore.scala 102:34]
  wire [1:0] frontend_io_out_0_bits_ctrl_src2Type; // @[NutCore.scala 102:34]
  wire [2:0] frontend_io_out_0_bits_ctrl_fuType; // @[NutCore.scala 102:34]
  wire [6:0] frontend_io_out_0_bits_ctrl_fuOpType; // @[NutCore.scala 102:34]
  wire [4:0] frontend_io_out_0_bits_ctrl_rfSrc1; // @[NutCore.scala 102:34]
  wire [4:0] frontend_io_out_0_bits_ctrl_rfSrc2; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_ctrl_rfWen; // @[NutCore.scala 102:34]
  wire [4:0] frontend_io_out_0_bits_ctrl_rfDest; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_ctrl_isNutCoreTrap; // @[NutCore.scala 102:34]
  wire [63:0] frontend_io_out_0_bits_data_imm; // @[NutCore.scala 102:34]
  wire  frontend_io_out_1_bits_cf_intrVec_0; // @[NutCore.scala 102:34]
  wire  frontend_io_out_1_bits_cf_intrVec_1; // @[NutCore.scala 102:34]
  wire  frontend_io_out_1_bits_cf_intrVec_2; // @[NutCore.scala 102:34]
  wire  frontend_io_out_1_bits_cf_intrVec_3; // @[NutCore.scala 102:34]
  wire  frontend_io_out_1_bits_cf_intrVec_4; // @[NutCore.scala 102:34]
  wire  frontend_io_out_1_bits_cf_intrVec_5; // @[NutCore.scala 102:34]
  wire  frontend_io_out_1_bits_cf_intrVec_6; // @[NutCore.scala 102:34]
  wire  frontend_io_out_1_bits_cf_intrVec_7; // @[NutCore.scala 102:34]
  wire  frontend_io_out_1_bits_cf_intrVec_8; // @[NutCore.scala 102:34]
  wire  frontend_io_out_1_bits_cf_intrVec_9; // @[NutCore.scala 102:34]
  wire  frontend_io_out_1_bits_cf_intrVec_10; // @[NutCore.scala 102:34]
  wire  frontend_io_out_1_bits_cf_intrVec_11; // @[NutCore.scala 102:34]
  wire  frontend_io_imem_req_ready; // @[NutCore.scala 102:34]
  wire  frontend_io_imem_req_valid; // @[NutCore.scala 102:34]
  wire [38:0] frontend_io_imem_req_bits_addr; // @[NutCore.scala 102:34]
  wire [86:0] frontend_io_imem_req_bits_user; // @[NutCore.scala 102:34]
  wire  frontend_io_imem_resp_ready; // @[NutCore.scala 102:34]
  wire  frontend_io_imem_resp_valid; // @[NutCore.scala 102:34]
  wire [63:0] frontend_io_imem_resp_bits_rdata; // @[NutCore.scala 102:34]
  wire [86:0] frontend_io_imem_resp_bits_user; // @[NutCore.scala 102:34]
  wire [3:0] frontend_io_flushVec; // @[NutCore.scala 102:34]
  wire  frontend_io_ipf; // @[NutCore.scala 102:34]
  wire [38:0] frontend_io_redirect_target; // @[NutCore.scala 102:34]
  wire  frontend_io_redirect_valid; // @[NutCore.scala 102:34]
  wire  frontend_flushICache; // @[NutCore.scala 102:34]
  wire  frontend__T_243_valid; // @[NutCore.scala 102:34]
  wire [38:0] frontend__T_243_pc; // @[NutCore.scala 102:34]
  wire  frontend__T_243_isMissPredict; // @[NutCore.scala 102:34]
  wire [38:0] frontend__T_243_actualTarget; // @[NutCore.scala 102:34]
  wire  frontend__T_243_actualTaken; // @[NutCore.scala 102:34]
  wire [6:0] frontend__T_243_fuOpType; // @[NutCore.scala 102:34]
  wire [1:0] frontend__T_243_btbType; // @[NutCore.scala 102:34]
  wire  frontend__T_243_isRVC; // @[NutCore.scala 102:34]
  wire  frontend_DISPLAY_ENABLE; // @[NutCore.scala 102:34]
  wire  frontend_vmEnable; // @[NutCore.scala 102:34]
  wire [11:0] frontend_intrVec; // @[NutCore.scala 102:34]
  wire  frontend__T_0; // @[NutCore.scala 102:34]
  wire  frontend__T_65; // @[NutCore.scala 102:34]
  wire  frontend_flushTLB; // @[NutCore.scala 102:34]
  wire  frontend__T_66; // @[NutCore.scala 102:34]
  wire  Backend_inorder_clock; // @[NutCore.scala 144:25]
  wire  Backend_inorder_reset; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_ready; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_valid; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder_io_in_0_bits_cf_instr; // @[NutCore.scala 144:25]
  wire [38:0] Backend_inorder_io_in_0_bits_cf_pc; // @[NutCore.scala 144:25]
  wire [38:0] Backend_inorder_io_in_0_bits_cf_pnpc; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_cf_exceptionVec_1; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_cf_exceptionVec_2; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_cf_exceptionVec_12; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_0; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_1; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_2; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_3; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_4; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_5; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_6; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_7; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_8; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_9; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_10; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_11; // @[NutCore.scala 144:25]
  wire [3:0] Backend_inorder_io_in_0_bits_cf_brIdx; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_cf_crossPageIPFFix; // @[NutCore.scala 144:25]
  wire [1:0] Backend_inorder_io_in_0_bits_ctrl_src1Type; // @[NutCore.scala 144:25]
  wire [1:0] Backend_inorder_io_in_0_bits_ctrl_src2Type; // @[NutCore.scala 144:25]
  wire [2:0] Backend_inorder_io_in_0_bits_ctrl_fuType; // @[NutCore.scala 144:25]
  wire [6:0] Backend_inorder_io_in_0_bits_ctrl_fuOpType; // @[NutCore.scala 144:25]
  wire [4:0] Backend_inorder_io_in_0_bits_ctrl_rfSrc1; // @[NutCore.scala 144:25]
  wire [4:0] Backend_inorder_io_in_0_bits_ctrl_rfSrc2; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_ctrl_rfWen; // @[NutCore.scala 144:25]
  wire [4:0] Backend_inorder_io_in_0_bits_ctrl_rfDest; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_ctrl_isNutCoreTrap; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder_io_in_0_bits_data_imm; // @[NutCore.scala 144:25]
  wire [1:0] Backend_inorder_io_flush; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_dmem_req_ready; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_dmem_req_valid; // @[NutCore.scala 144:25]
  wire [38:0] Backend_inorder_io_dmem_req_bits_addr; // @[NutCore.scala 144:25]
  wire [2:0] Backend_inorder_io_dmem_req_bits_size; // @[NutCore.scala 144:25]
  wire [3:0] Backend_inorder_io_dmem_req_bits_cmd; // @[NutCore.scala 144:25]
  wire [7:0] Backend_inorder_io_dmem_req_bits_wmask; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder_io_dmem_req_bits_wdata; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_dmem_resp_valid; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder_io_dmem_resp_bits_rdata; // @[NutCore.scala 144:25]
  wire [1:0] Backend_inorder_io_memMMU_imem_priviledgeMode; // @[NutCore.scala 144:25]
  wire [1:0] Backend_inorder_io_memMMU_dmem_priviledgeMode; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_memMMU_dmem_status_sum; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_memMMU_dmem_status_mxr; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_memMMU_dmem_loadPF; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_memMMU_dmem_storePF; // @[NutCore.scala 144:25]
  wire [38:0] Backend_inorder_io_memMMU_dmem_addr; // @[NutCore.scala 144:25]
  wire [38:0] Backend_inorder_io_redirect_target; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_redirect_valid; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_4181; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_4184; // @[NutCore.scala 144:25]
  wire  Backend_inorder__T_38; // @[NutCore.scala 144:25]
  wire  Backend_inorder_flushICache; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_4185; // @[NutCore.scala 144:25]
  wire  Backend_inorder_falseWire; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder_satp; // @[NutCore.scala 144:25]
  wire  Backend_inorder__T_243_valid; // @[NutCore.scala 144:25]
  wire [38:0] Backend_inorder__T_243_pc; // @[NutCore.scala 144:25]
  wire  Backend_inorder__T_243_isMissPredict; // @[NutCore.scala 144:25]
  wire [38:0] Backend_inorder__T_243_actualTarget; // @[NutCore.scala 144:25]
  wire  Backend_inorder__T_243_actualTaken; // @[NutCore.scala 144:25]
  wire [6:0] Backend_inorder__T_243_fuOpType; // @[NutCore.scala 144:25]
  wire [1:0] Backend_inorder__T_243_btbType; // @[NutCore.scala 144:25]
  wire  Backend_inorder__T_243_isRVC; // @[NutCore.scala 144:25]
  wire  Backend_inorder_falseWire_0; // @[NutCore.scala 144:25]
  wire [1:0] Backend_inorder__T_4178; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_284_0; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_284_1; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_284_2; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_284_3; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_284_4; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_284_5; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_284_6; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_284_7; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_284_8; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_284_9; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_284_10; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_284_11; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_284_12; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_284_13; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_284_14; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_284_15; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_284_16; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_284_17; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_284_18; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_284_19; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_284_20; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_284_21; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_284_22; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_284_23; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_284_24; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_284_25; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_284_26; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_284_27; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_284_28; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_284_29; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_284_30; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_284_31; // @[NutCore.scala 144:25]
  wire  Backend_inorder_mmio; // @[NutCore.scala 144:25]
  wire  Backend_inorder__T_36; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_extra_mtip; // @[NutCore.scala 144:25]
  wire  Backend_inorder_amoReq; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_32; // @[NutCore.scala 144:25]
  wire  Backend_inorder__T_13; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_extra_meip_0; // @[NutCore.scala 144:25]
  wire  Backend_inorder_vmEnable; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_31; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_37; // @[NutCore.scala 144:25]
  wire  Backend_inorder__T_26; // @[NutCore.scala 144:25]
  wire [11:0] Backend_inorder_intrVec; // @[NutCore.scala 144:25]
  wire  Backend_inorder__T_37_0; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_extra_msip; // @[NutCore.scala 144:25]
  wire  Backend_inorder__T_65; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_4183; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_4182; // @[NutCore.scala 144:25]
  wire  Backend_inorder_flushTLB; // @[NutCore.scala 144:25]
  wire  Backend_inorder__T_33; // @[NutCore.scala 144:25]
  wire  Backend_inorder__T_66; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder__T_4179; // @[NutCore.scala 144:25]
  wire  SimpleBusCrossbarNto1_clock; // @[NutCore.scala 148:26]
  wire  SimpleBusCrossbarNto1_reset; // @[NutCore.scala 148:26]
  wire  SimpleBusCrossbarNto1_io_in_0_req_ready; // @[NutCore.scala 148:26]
  wire  SimpleBusCrossbarNto1_io_in_0_req_valid; // @[NutCore.scala 148:26]
  wire [31:0] SimpleBusCrossbarNto1_io_in_0_req_bits_addr; // @[NutCore.scala 148:26]
  wire [3:0] SimpleBusCrossbarNto1_io_in_0_req_bits_cmd; // @[NutCore.scala 148:26]
  wire [7:0] SimpleBusCrossbarNto1_io_in_0_req_bits_wmask; // @[NutCore.scala 148:26]
  wire [63:0] SimpleBusCrossbarNto1_io_in_0_req_bits_wdata; // @[NutCore.scala 148:26]
  wire  SimpleBusCrossbarNto1_io_in_0_resp_valid; // @[NutCore.scala 148:26]
  wire [3:0] SimpleBusCrossbarNto1_io_in_0_resp_bits_cmd; // @[NutCore.scala 148:26]
  wire [63:0] SimpleBusCrossbarNto1_io_in_0_resp_bits_rdata; // @[NutCore.scala 148:26]
  wire  SimpleBusCrossbarNto1_io_in_1_req_ready; // @[NutCore.scala 148:26]
  wire  SimpleBusCrossbarNto1_io_in_1_req_valid; // @[NutCore.scala 148:26]
  wire [31:0] SimpleBusCrossbarNto1_io_in_1_req_bits_addr; // @[NutCore.scala 148:26]
  wire [2:0] SimpleBusCrossbarNto1_io_in_1_req_bits_size; // @[NutCore.scala 148:26]
  wire [3:0] SimpleBusCrossbarNto1_io_in_1_req_bits_cmd; // @[NutCore.scala 148:26]
  wire [7:0] SimpleBusCrossbarNto1_io_in_1_req_bits_wmask; // @[NutCore.scala 148:26]
  wire [63:0] SimpleBusCrossbarNto1_io_in_1_req_bits_wdata; // @[NutCore.scala 148:26]
  wire  SimpleBusCrossbarNto1_io_in_1_resp_valid; // @[NutCore.scala 148:26]
  wire [3:0] SimpleBusCrossbarNto1_io_in_1_resp_bits_cmd; // @[NutCore.scala 148:26]
  wire [63:0] SimpleBusCrossbarNto1_io_in_1_resp_bits_rdata; // @[NutCore.scala 148:26]
  wire  SimpleBusCrossbarNto1_io_out_req_ready; // @[NutCore.scala 148:26]
  wire  SimpleBusCrossbarNto1_io_out_req_valid; // @[NutCore.scala 148:26]
  wire [31:0] SimpleBusCrossbarNto1_io_out_req_bits_addr; // @[NutCore.scala 148:26]
  wire [2:0] SimpleBusCrossbarNto1_io_out_req_bits_size; // @[NutCore.scala 148:26]
  wire [3:0] SimpleBusCrossbarNto1_io_out_req_bits_cmd; // @[NutCore.scala 148:26]
  wire [7:0] SimpleBusCrossbarNto1_io_out_req_bits_wmask; // @[NutCore.scala 148:26]
  wire [63:0] SimpleBusCrossbarNto1_io_out_req_bits_wdata; // @[NutCore.scala 148:26]
  wire  SimpleBusCrossbarNto1_io_out_resp_ready; // @[NutCore.scala 148:26]
  wire  SimpleBusCrossbarNto1_io_out_resp_valid; // @[NutCore.scala 148:26]
  wire [3:0] SimpleBusCrossbarNto1_io_out_resp_bits_cmd; // @[NutCore.scala 148:26]
  wire [63:0] SimpleBusCrossbarNto1_io_out_resp_bits_rdata; // @[NutCore.scala 148:26]
  wire  SimpleBusCrossbarNto1_1_clock; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_reset; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_in_0_req_ready; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_in_0_req_valid; // @[NutCore.scala 149:26]
  wire [31:0] SimpleBusCrossbarNto1_1_io_in_0_req_bits_addr; // @[NutCore.scala 149:26]
  wire [2:0] SimpleBusCrossbarNto1_1_io_in_0_req_bits_size; // @[NutCore.scala 149:26]
  wire [3:0] SimpleBusCrossbarNto1_1_io_in_0_req_bits_cmd; // @[NutCore.scala 149:26]
  wire [7:0] SimpleBusCrossbarNto1_1_io_in_0_req_bits_wmask; // @[NutCore.scala 149:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_in_0_req_bits_wdata; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_in_0_resp_valid; // @[NutCore.scala 149:26]
  wire [3:0] SimpleBusCrossbarNto1_1_io_in_0_resp_bits_cmd; // @[NutCore.scala 149:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_in_0_resp_bits_rdata; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_in_1_req_ready; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_in_1_req_valid; // @[NutCore.scala 149:26]
  wire [31:0] SimpleBusCrossbarNto1_1_io_in_1_req_bits_addr; // @[NutCore.scala 149:26]
  wire [3:0] SimpleBusCrossbarNto1_1_io_in_1_req_bits_cmd; // @[NutCore.scala 149:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_in_1_req_bits_wdata; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_in_1_resp_valid; // @[NutCore.scala 149:26]
  wire [3:0] SimpleBusCrossbarNto1_1_io_in_1_resp_bits_cmd; // @[NutCore.scala 149:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_in_1_resp_bits_rdata; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_in_2_req_ready; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_in_2_req_valid; // @[NutCore.scala 149:26]
  wire [31:0] SimpleBusCrossbarNto1_1_io_in_2_req_bits_addr; // @[NutCore.scala 149:26]
  wire [3:0] SimpleBusCrossbarNto1_1_io_in_2_req_bits_cmd; // @[NutCore.scala 149:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_in_2_req_bits_wdata; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_in_2_resp_valid; // @[NutCore.scala 149:26]
  wire [3:0] SimpleBusCrossbarNto1_1_io_in_2_resp_bits_cmd; // @[NutCore.scala 149:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_in_2_resp_bits_rdata; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_in_3_req_ready; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_in_3_req_valid; // @[NutCore.scala 149:26]
  wire [31:0] SimpleBusCrossbarNto1_1_io_in_3_req_bits_addr; // @[NutCore.scala 149:26]
  wire [2:0] SimpleBusCrossbarNto1_1_io_in_3_req_bits_size; // @[NutCore.scala 149:26]
  wire [3:0] SimpleBusCrossbarNto1_1_io_in_3_req_bits_cmd; // @[NutCore.scala 149:26]
  wire [7:0] SimpleBusCrossbarNto1_1_io_in_3_req_bits_wmask; // @[NutCore.scala 149:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_in_3_req_bits_wdata; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_in_3_resp_ready; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_in_3_resp_valid; // @[NutCore.scala 149:26]
  wire [3:0] SimpleBusCrossbarNto1_1_io_in_3_resp_bits_cmd; // @[NutCore.scala 149:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_in_3_resp_bits_rdata; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_out_req_ready; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_out_req_valid; // @[NutCore.scala 149:26]
  wire [31:0] SimpleBusCrossbarNto1_1_io_out_req_bits_addr; // @[NutCore.scala 149:26]
  wire [2:0] SimpleBusCrossbarNto1_1_io_out_req_bits_size; // @[NutCore.scala 149:26]
  wire [3:0] SimpleBusCrossbarNto1_1_io_out_req_bits_cmd; // @[NutCore.scala 149:26]
  wire [7:0] SimpleBusCrossbarNto1_1_io_out_req_bits_wmask; // @[NutCore.scala 149:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_out_req_bits_wdata; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_out_resp_ready; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_out_resp_valid; // @[NutCore.scala 149:26]
  wire [3:0] SimpleBusCrossbarNto1_1_io_out_resp_bits_cmd; // @[NutCore.scala 149:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_out_resp_bits_rdata; // @[NutCore.scala 149:26]
  wire  EmbeddedTLB_clock; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_reset; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_in_req_ready; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_in_req_valid; // @[EmbeddedTLB.scala 427:23]
  wire [38:0] EmbeddedTLB_io_in_req_bits_addr; // @[EmbeddedTLB.scala 427:23]
  wire [86:0] EmbeddedTLB_io_in_req_bits_user; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_in_resp_ready; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_in_resp_valid; // @[EmbeddedTLB.scala 427:23]
  wire [3:0] EmbeddedTLB_io_in_resp_bits_cmd; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_io_in_resp_bits_rdata; // @[EmbeddedTLB.scala 427:23]
  wire [86:0] EmbeddedTLB_io_in_resp_bits_user; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_out_req_ready; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_out_req_valid; // @[EmbeddedTLB.scala 427:23]
  wire [31:0] EmbeddedTLB_io_out_req_bits_addr; // @[EmbeddedTLB.scala 427:23]
  wire [3:0] EmbeddedTLB_io_out_req_bits_cmd; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_io_out_req_bits_wdata; // @[EmbeddedTLB.scala 427:23]
  wire [86:0] EmbeddedTLB_io_out_req_bits_user; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_out_resp_ready; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_out_resp_valid; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_io_out_resp_bits_rdata; // @[EmbeddedTLB.scala 427:23]
  wire [86:0] EmbeddedTLB_io_out_resp_bits_user; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_mem_req_ready; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_mem_req_valid; // @[EmbeddedTLB.scala 427:23]
  wire [31:0] EmbeddedTLB_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 427:23]
  wire [3:0] EmbeddedTLB_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_mem_resp_valid; // @[EmbeddedTLB.scala 427:23]
  wire [3:0] EmbeddedTLB_io_mem_resp_bits_cmd; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_io_mem_resp_bits_rdata; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_flush; // @[EmbeddedTLB.scala 427:23]
  wire [1:0] EmbeddedTLB_io_csrMMU_priviledgeMode; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_csrMMU_loadPF; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_csrMMU_storePF; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_cacheEmpty; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_ipf; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_CSRSATP; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_DISPLAY_ENABLE; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_MOUFlushTLB; // @[EmbeddedTLB.scala 427:23]
  wire  Cache_clock; // @[Cache.scala 678:35]
  wire  Cache_reset; // @[Cache.scala 678:35]
  wire  Cache_io_in_req_ready; // @[Cache.scala 678:35]
  wire  Cache_io_in_req_valid; // @[Cache.scala 678:35]
  wire [31:0] Cache_io_in_req_bits_addr; // @[Cache.scala 678:35]
  wire [86:0] Cache_io_in_req_bits_user; // @[Cache.scala 678:35]
  wire  Cache_io_in_resp_ready; // @[Cache.scala 678:35]
  wire  Cache_io_in_resp_valid; // @[Cache.scala 678:35]
  wire [63:0] Cache_io_in_resp_bits_rdata; // @[Cache.scala 678:35]
  wire [86:0] Cache_io_in_resp_bits_user; // @[Cache.scala 678:35]
  wire [1:0] Cache_io_flush; // @[Cache.scala 678:35]
  wire  Cache_io_out_mem_req_ready; // @[Cache.scala 678:35]
  wire  Cache_io_out_mem_req_valid; // @[Cache.scala 678:35]
  wire [31:0] Cache_io_out_mem_req_bits_addr; // @[Cache.scala 678:35]
  wire [3:0] Cache_io_out_mem_req_bits_cmd; // @[Cache.scala 678:35]
  wire [63:0] Cache_io_out_mem_req_bits_wdata; // @[Cache.scala 678:35]
  wire  Cache_io_out_mem_resp_valid; // @[Cache.scala 678:35]
  wire [3:0] Cache_io_out_mem_resp_bits_cmd; // @[Cache.scala 678:35]
  wire [63:0] Cache_io_out_mem_resp_bits_rdata; // @[Cache.scala 678:35]
  wire  Cache_io_mmio_req_ready; // @[Cache.scala 678:35]
  wire  Cache_io_mmio_req_valid; // @[Cache.scala 678:35]
  wire [31:0] Cache_io_mmio_req_bits_addr; // @[Cache.scala 678:35]
  wire  Cache_io_mmio_resp_valid; // @[Cache.scala 678:35]
  wire [63:0] Cache_io_mmio_resp_bits_rdata; // @[Cache.scala 678:35]
  wire  Cache_io_empty; // @[Cache.scala 678:35]
  wire  Cache_MOUFlushICache; // @[Cache.scala 678:35]
  wire  Cache_DISPLAY_ENABLE; // @[Cache.scala 678:35]
  wire  EmbeddedTLB_1_clock; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_reset; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_in_req_ready; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_in_req_valid; // @[EmbeddedTLB.scala 427:23]
  wire [38:0] EmbeddedTLB_1_io_in_req_bits_addr; // @[EmbeddedTLB.scala 427:23]
  wire [2:0] EmbeddedTLB_1_io_in_req_bits_size; // @[EmbeddedTLB.scala 427:23]
  wire [3:0] EmbeddedTLB_1_io_in_req_bits_cmd; // @[EmbeddedTLB.scala 427:23]
  wire [7:0] EmbeddedTLB_1_io_in_req_bits_wmask; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_1_io_in_req_bits_wdata; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_in_resp_valid; // @[EmbeddedTLB.scala 427:23]
  wire [3:0] EmbeddedTLB_1_io_in_resp_bits_cmd; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_1_io_in_resp_bits_rdata; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_out_req_ready; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_out_req_valid; // @[EmbeddedTLB.scala 427:23]
  wire [31:0] EmbeddedTLB_1_io_out_req_bits_addr; // @[EmbeddedTLB.scala 427:23]
  wire [2:0] EmbeddedTLB_1_io_out_req_bits_size; // @[EmbeddedTLB.scala 427:23]
  wire [3:0] EmbeddedTLB_1_io_out_req_bits_cmd; // @[EmbeddedTLB.scala 427:23]
  wire [7:0] EmbeddedTLB_1_io_out_req_bits_wmask; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_1_io_out_req_bits_wdata; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_out_resp_ready; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_out_resp_valid; // @[EmbeddedTLB.scala 427:23]
  wire [3:0] EmbeddedTLB_1_io_out_resp_bits_cmd; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_1_io_out_resp_bits_rdata; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_mem_req_ready; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_mem_req_valid; // @[EmbeddedTLB.scala 427:23]
  wire [31:0] EmbeddedTLB_1_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 427:23]
  wire [3:0] EmbeddedTLB_1_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_1_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_mem_resp_valid; // @[EmbeddedTLB.scala 427:23]
  wire [3:0] EmbeddedTLB_1_io_mem_resp_bits_cmd; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_1_io_mem_resp_bits_rdata; // @[EmbeddedTLB.scala 427:23]
  wire [1:0] EmbeddedTLB_1_io_csrMMU_priviledgeMode; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_csrMMU_status_sum; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_csrMMU_status_mxr; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_csrMMU_loadPF; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_csrMMU_storePF; // @[EmbeddedTLB.scala 427:23]
  wire [38:0] EmbeddedTLB_1_io_csrMMU_addr; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_cacheEmpty; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_ipf; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1__T_38_0; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_1_CSRSATP; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_amoReq; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_DISPLAY_ENABLE; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_vmEnable_0; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1__T_37_1; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_MOUFlushTLB; // @[EmbeddedTLB.scala 427:23]
  wire  Cache_1_clock; // @[Cache.scala 678:35]
  wire  Cache_1_reset; // @[Cache.scala 678:35]
  wire  Cache_1_io_in_req_ready; // @[Cache.scala 678:35]
  wire  Cache_1_io_in_req_valid; // @[Cache.scala 678:35]
  wire [31:0] Cache_1_io_in_req_bits_addr; // @[Cache.scala 678:35]
  wire [2:0] Cache_1_io_in_req_bits_size; // @[Cache.scala 678:35]
  wire [3:0] Cache_1_io_in_req_bits_cmd; // @[Cache.scala 678:35]
  wire [7:0] Cache_1_io_in_req_bits_wmask; // @[Cache.scala 678:35]
  wire [63:0] Cache_1_io_in_req_bits_wdata; // @[Cache.scala 678:35]
  wire  Cache_1_io_in_resp_ready; // @[Cache.scala 678:35]
  wire  Cache_1_io_in_resp_valid; // @[Cache.scala 678:35]
  wire [3:0] Cache_1_io_in_resp_bits_cmd; // @[Cache.scala 678:35]
  wire [63:0] Cache_1_io_in_resp_bits_rdata; // @[Cache.scala 678:35]
  wire  Cache_1_io_out_mem_req_ready; // @[Cache.scala 678:35]
  wire  Cache_1_io_out_mem_req_valid; // @[Cache.scala 678:35]
  wire [31:0] Cache_1_io_out_mem_req_bits_addr; // @[Cache.scala 678:35]
  wire [3:0] Cache_1_io_out_mem_req_bits_cmd; // @[Cache.scala 678:35]
  wire [63:0] Cache_1_io_out_mem_req_bits_wdata; // @[Cache.scala 678:35]
  wire  Cache_1_io_out_mem_resp_valid; // @[Cache.scala 678:35]
  wire [3:0] Cache_1_io_out_mem_resp_bits_cmd; // @[Cache.scala 678:35]
  wire [63:0] Cache_1_io_out_mem_resp_bits_rdata; // @[Cache.scala 678:35]
  wire  Cache_1_io_out_coh_req_ready; // @[Cache.scala 678:35]
  wire  Cache_1_io_out_coh_req_valid; // @[Cache.scala 678:35]
  wire [31:0] Cache_1_io_out_coh_req_bits_addr; // @[Cache.scala 678:35]
  wire [63:0] Cache_1_io_out_coh_req_bits_wdata; // @[Cache.scala 678:35]
  wire  Cache_1_io_out_coh_resp_valid; // @[Cache.scala 678:35]
  wire [3:0] Cache_1_io_out_coh_resp_bits_cmd; // @[Cache.scala 678:35]
  wire [63:0] Cache_1_io_out_coh_resp_bits_rdata; // @[Cache.scala 678:35]
  wire  Cache_1_io_mmio_req_ready; // @[Cache.scala 678:35]
  wire  Cache_1_io_mmio_req_valid; // @[Cache.scala 678:35]
  wire [31:0] Cache_1_io_mmio_req_bits_addr; // @[Cache.scala 678:35]
  wire [2:0] Cache_1_io_mmio_req_bits_size; // @[Cache.scala 678:35]
  wire [3:0] Cache_1_io_mmio_req_bits_cmd; // @[Cache.scala 678:35]
  wire [7:0] Cache_1_io_mmio_req_bits_wmask; // @[Cache.scala 678:35]
  wire [63:0] Cache_1_io_mmio_req_bits_wdata; // @[Cache.scala 678:35]
  wire  Cache_1_io_mmio_resp_valid; // @[Cache.scala 678:35]
  wire [63:0] Cache_1_io_mmio_resp_bits_rdata; // @[Cache.scala 678:35]
  wire  Cache_1_io_empty; // @[Cache.scala 678:35]
  wire  Cache_1_mmio; // @[Cache.scala 678:35]
  wire  Cache_1_DISPLAY_ENABLE; // @[Cache.scala 678:35]
  reg [63:0] _T_6_0_cf_instr; // @[PipelineVector.scala 29:29]
  reg [38:0] _T_6_0_cf_pc; // @[PipelineVector.scala 29:29]
  reg [38:0] _T_6_0_cf_pnpc; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_cf_exceptionVec_1; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_cf_exceptionVec_2; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_cf_exceptionVec_12; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_cf_intrVec_0; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_cf_intrVec_1; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_cf_intrVec_2; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_cf_intrVec_3; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_cf_intrVec_4; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_cf_intrVec_5; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_cf_intrVec_6; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_cf_intrVec_7; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_cf_intrVec_8; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_cf_intrVec_9; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_cf_intrVec_10; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_cf_intrVec_11; // @[PipelineVector.scala 29:29]
  reg [3:0] _T_6_0_cf_brIdx; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29]
  reg [1:0] _T_6_0_ctrl_src1Type; // @[PipelineVector.scala 29:29]
  reg [1:0] _T_6_0_ctrl_src2Type; // @[PipelineVector.scala 29:29]
  reg [2:0] _T_6_0_ctrl_fuType; // @[PipelineVector.scala 29:29]
  reg [6:0] _T_6_0_ctrl_fuOpType; // @[PipelineVector.scala 29:29]
  reg [4:0] _T_6_0_ctrl_rfSrc1; // @[PipelineVector.scala 29:29]
  reg [4:0] _T_6_0_ctrl_rfSrc2; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_ctrl_rfWen; // @[PipelineVector.scala 29:29]
  reg [4:0] _T_6_0_ctrl_rfDest; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_ctrl_isNutCoreTrap; // @[PipelineVector.scala 29:29]
  reg [63:0] _T_6_0_data_imm; // @[PipelineVector.scala 29:29]
  reg [63:0] _T_6_1_cf_instr; // @[PipelineVector.scala 29:29]
  reg [38:0] _T_6_1_cf_pc; // @[PipelineVector.scala 29:29]
  reg [38:0] _T_6_1_cf_pnpc; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_cf_exceptionVec_1; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_cf_exceptionVec_2; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_cf_exceptionVec_12; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_cf_intrVec_0; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_cf_intrVec_1; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_cf_intrVec_2; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_cf_intrVec_3; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_cf_intrVec_4; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_cf_intrVec_5; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_cf_intrVec_6; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_cf_intrVec_7; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_cf_intrVec_8; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_cf_intrVec_9; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_cf_intrVec_10; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_cf_intrVec_11; // @[PipelineVector.scala 29:29]
  reg [3:0] _T_6_1_cf_brIdx; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29]
  reg [1:0] _T_6_1_ctrl_src1Type; // @[PipelineVector.scala 29:29]
  reg [1:0] _T_6_1_ctrl_src2Type; // @[PipelineVector.scala 29:29]
  reg [2:0] _T_6_1_ctrl_fuType; // @[PipelineVector.scala 29:29]
  reg [6:0] _T_6_1_ctrl_fuOpType; // @[PipelineVector.scala 29:29]
  reg [4:0] _T_6_1_ctrl_rfSrc1; // @[PipelineVector.scala 29:29]
  reg [4:0] _T_6_1_ctrl_rfSrc2; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_ctrl_rfWen; // @[PipelineVector.scala 29:29]
  reg [4:0] _T_6_1_ctrl_rfDest; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_ctrl_isNutCoreTrap; // @[PipelineVector.scala 29:29]
  reg [63:0] _T_6_1_data_imm; // @[PipelineVector.scala 29:29]
  reg [63:0] _T_6_2_cf_instr; // @[PipelineVector.scala 29:29]
  reg [38:0] _T_6_2_cf_pc; // @[PipelineVector.scala 29:29]
  reg [38:0] _T_6_2_cf_pnpc; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_cf_exceptionVec_1; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_cf_exceptionVec_2; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_cf_exceptionVec_12; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_cf_intrVec_0; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_cf_intrVec_1; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_cf_intrVec_2; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_cf_intrVec_3; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_cf_intrVec_4; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_cf_intrVec_5; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_cf_intrVec_6; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_cf_intrVec_7; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_cf_intrVec_8; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_cf_intrVec_9; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_cf_intrVec_10; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_cf_intrVec_11; // @[PipelineVector.scala 29:29]
  reg [3:0] _T_6_2_cf_brIdx; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29]
  reg [1:0] _T_6_2_ctrl_src1Type; // @[PipelineVector.scala 29:29]
  reg [1:0] _T_6_2_ctrl_src2Type; // @[PipelineVector.scala 29:29]
  reg [2:0] _T_6_2_ctrl_fuType; // @[PipelineVector.scala 29:29]
  reg [6:0] _T_6_2_ctrl_fuOpType; // @[PipelineVector.scala 29:29]
  reg [4:0] _T_6_2_ctrl_rfSrc1; // @[PipelineVector.scala 29:29]
  reg [4:0] _T_6_2_ctrl_rfSrc2; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_ctrl_rfWen; // @[PipelineVector.scala 29:29]
  reg [4:0] _T_6_2_ctrl_rfDest; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_ctrl_isNutCoreTrap; // @[PipelineVector.scala 29:29]
  reg [63:0] _T_6_2_data_imm; // @[PipelineVector.scala 29:29]
  reg [63:0] _T_6_3_cf_instr; // @[PipelineVector.scala 29:29]
  reg [38:0] _T_6_3_cf_pc; // @[PipelineVector.scala 29:29]
  reg [38:0] _T_6_3_cf_pnpc; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_cf_exceptionVec_1; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_cf_exceptionVec_2; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_cf_exceptionVec_12; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_cf_intrVec_0; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_cf_intrVec_1; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_cf_intrVec_2; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_cf_intrVec_3; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_cf_intrVec_4; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_cf_intrVec_5; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_cf_intrVec_6; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_cf_intrVec_7; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_cf_intrVec_8; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_cf_intrVec_9; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_cf_intrVec_10; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_cf_intrVec_11; // @[PipelineVector.scala 29:29]
  reg [3:0] _T_6_3_cf_brIdx; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29]
  reg [1:0] _T_6_3_ctrl_src1Type; // @[PipelineVector.scala 29:29]
  reg [1:0] _T_6_3_ctrl_src2Type; // @[PipelineVector.scala 29:29]
  reg [2:0] _T_6_3_ctrl_fuType; // @[PipelineVector.scala 29:29]
  reg [6:0] _T_6_3_ctrl_fuOpType; // @[PipelineVector.scala 29:29]
  reg [4:0] _T_6_3_ctrl_rfSrc1; // @[PipelineVector.scala 29:29]
  reg [4:0] _T_6_3_ctrl_rfSrc2; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_ctrl_rfWen; // @[PipelineVector.scala 29:29]
  reg [4:0] _T_6_3_ctrl_rfDest; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_ctrl_isNutCoreTrap; // @[PipelineVector.scala 29:29]
  reg [63:0] _T_6_3_data_imm; // @[PipelineVector.scala 29:29]
  reg [1:0] _T_7; // @[PipelineVector.scala 30:33]
  reg [1:0] _T_8; // @[PipelineVector.scala 31:33]
  wire [1:0] _T_11 = _T_7 + 2'h1; // @[PipelineVector.scala 33:63]
  wire  _T_12 = _T_11 != _T_8; // @[PipelineVector.scala 33:74]
  wire [1:0] _T_14 = _T_7 + 2'h2; // @[PipelineVector.scala 33:63]
  wire  _T_15 = _T_14 != _T_8; // @[PipelineVector.scala 33:74]
  wire  _T_17 = _T_12 & _T_15; // @[PipelineVector.scala 33:124]
  wire  _T_18_0 = frontend_io_out_0_valid; // @[PipelineVector.scala 36:27 PipelineVector.scala 37:20]
  wire [1:0] _T_19 = {{1'd0}, _T_18_0}; // @[PipelineVector.scala 40:46]
  wire  _T_20 = _T_19 >= 2'h1; // @[PipelineVector.scala 41:53]
  wire  _T_21 = _T_19 >= 2'h2; // @[PipelineVector.scala 41:53]
  wire  _T_22 = frontend_io_out_0_ready & frontend_io_out_0_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _T_25 = {{1'd0}, _T_7}; // @[PipelineVector.scala 45:45]
  wire [63:0] _T_27_cf_instr = _T_18_0 ? frontend_io_out_0_bits_cf_instr : 64'h0; // @[PipelineVector.scala 45:69]
  wire [38:0] _T_27_cf_pc = _T_18_0 ? frontend_io_out_0_bits_cf_pc : 39'h0; // @[PipelineVector.scala 45:69]
  wire [38:0] _T_27_cf_pnpc = _T_18_0 ? frontend_io_out_0_bits_cf_pnpc : 39'h0; // @[PipelineVector.scala 45:69]
  wire  _T_27_cf_exceptionVec_1 = _T_18_0 & frontend_io_out_0_bits_cf_exceptionVec_1; // @[PipelineVector.scala 45:69]
  wire  _T_27_cf_exceptionVec_2 = _T_18_0 & frontend_io_out_0_bits_cf_exceptionVec_2; // @[PipelineVector.scala 45:69]
  wire  _T_27_cf_exceptionVec_12 = _T_18_0 & frontend_io_out_0_bits_cf_exceptionVec_12; // @[PipelineVector.scala 45:69]
  wire  _T_27_cf_intrVec_0 = _T_18_0 ? frontend_io_out_0_bits_cf_intrVec_0 : frontend_io_out_1_bits_cf_intrVec_0; // @[PipelineVector.scala 45:69]
  wire  _T_27_cf_intrVec_1 = _T_18_0 ? frontend_io_out_0_bits_cf_intrVec_1 : frontend_io_out_1_bits_cf_intrVec_1; // @[PipelineVector.scala 45:69]
  wire  _T_27_cf_intrVec_2 = _T_18_0 ? frontend_io_out_0_bits_cf_intrVec_2 : frontend_io_out_1_bits_cf_intrVec_2; // @[PipelineVector.scala 45:69]
  wire  _T_27_cf_intrVec_3 = _T_18_0 ? frontend_io_out_0_bits_cf_intrVec_3 : frontend_io_out_1_bits_cf_intrVec_3; // @[PipelineVector.scala 45:69]
  wire  _T_27_cf_intrVec_4 = _T_18_0 ? frontend_io_out_0_bits_cf_intrVec_4 : frontend_io_out_1_bits_cf_intrVec_4; // @[PipelineVector.scala 45:69]
  wire  _T_27_cf_intrVec_5 = _T_18_0 ? frontend_io_out_0_bits_cf_intrVec_5 : frontend_io_out_1_bits_cf_intrVec_5; // @[PipelineVector.scala 45:69]
  wire  _T_27_cf_intrVec_6 = _T_18_0 ? frontend_io_out_0_bits_cf_intrVec_6 : frontend_io_out_1_bits_cf_intrVec_6; // @[PipelineVector.scala 45:69]
  wire  _T_27_cf_intrVec_7 = _T_18_0 ? frontend_io_out_0_bits_cf_intrVec_7 : frontend_io_out_1_bits_cf_intrVec_7; // @[PipelineVector.scala 45:69]
  wire  _T_27_cf_intrVec_8 = _T_18_0 ? frontend_io_out_0_bits_cf_intrVec_8 : frontend_io_out_1_bits_cf_intrVec_8; // @[PipelineVector.scala 45:69]
  wire  _T_27_cf_intrVec_9 = _T_18_0 ? frontend_io_out_0_bits_cf_intrVec_9 : frontend_io_out_1_bits_cf_intrVec_9; // @[PipelineVector.scala 45:69]
  wire  _T_27_cf_intrVec_10 = _T_18_0 ? frontend_io_out_0_bits_cf_intrVec_10 : frontend_io_out_1_bits_cf_intrVec_10; // @[PipelineVector.scala 45:69]
  wire  _T_27_cf_intrVec_11 = _T_18_0 ? frontend_io_out_0_bits_cf_intrVec_11 : frontend_io_out_1_bits_cf_intrVec_11; // @[PipelineVector.scala 45:69]
  wire [3:0] _T_27_cf_brIdx = _T_18_0 ? frontend_io_out_0_bits_cf_brIdx : 4'h0; // @[PipelineVector.scala 45:69]
  wire  _T_27_cf_crossPageIPFFix = _T_18_0 & frontend_io_out_0_bits_cf_crossPageIPFFix; // @[PipelineVector.scala 45:69]
  wire [1:0] _T_27_ctrl_src1Type = _T_18_0 ? frontend_io_out_0_bits_ctrl_src1Type : 2'h1; // @[PipelineVector.scala 45:69]
  wire [1:0] _T_27_ctrl_src2Type = _T_18_0 ? frontend_io_out_0_bits_ctrl_src2Type : 2'h1; // @[PipelineVector.scala 45:69]
  wire [2:0] _T_27_ctrl_fuType = _T_18_0 ? frontend_io_out_0_bits_ctrl_fuType : 3'h3; // @[PipelineVector.scala 45:69]
  wire [6:0] _T_27_ctrl_fuOpType = _T_18_0 ? frontend_io_out_0_bits_ctrl_fuOpType : 7'h0; // @[PipelineVector.scala 45:69]
  wire [4:0] _T_27_ctrl_rfSrc1 = _T_18_0 ? frontend_io_out_0_bits_ctrl_rfSrc1 : 5'h0; // @[PipelineVector.scala 45:69]
  wire [4:0] _T_27_ctrl_rfSrc2 = _T_18_0 ? frontend_io_out_0_bits_ctrl_rfSrc2 : 5'h0; // @[PipelineVector.scala 45:69]
  wire  _T_27_ctrl_rfWen = _T_18_0 & frontend_io_out_0_bits_ctrl_rfWen; // @[PipelineVector.scala 45:69]
  wire [4:0] _T_27_ctrl_rfDest = _T_18_0 ? frontend_io_out_0_bits_ctrl_rfDest : 5'h0; // @[PipelineVector.scala 45:69]
  wire  _T_27_ctrl_isNutCoreTrap = _T_18_0 & frontend_io_out_0_bits_ctrl_isNutCoreTrap; // @[PipelineVector.scala 45:69]
  wire [63:0] _T_27_data_imm = _T_18_0 ? frontend_io_out_0_bits_data_imm : 64'h0; // @[PipelineVector.scala 45:69]
  wire [1:0] _T_29 = 2'h1 + _T_7; // @[PipelineVector.scala 46:45]
  wire  _T_6_T_29_cf_intrVec_0 = frontend_io_out_1_bits_cf_intrVec_0; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire  _T_6_T_29_cf_intrVec_1 = frontend_io_out_1_bits_cf_intrVec_1; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire  _T_6_T_29_cf_intrVec_2 = frontend_io_out_1_bits_cf_intrVec_2; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire  _T_6_T_29_cf_intrVec_3 = frontend_io_out_1_bits_cf_intrVec_3; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire  _T_6_T_29_cf_intrVec_4 = frontend_io_out_1_bits_cf_intrVec_4; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire  _T_6_T_29_cf_intrVec_5 = frontend_io_out_1_bits_cf_intrVec_5; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire  _T_6_T_29_cf_intrVec_6 = frontend_io_out_1_bits_cf_intrVec_6; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire  _T_6_T_29_cf_intrVec_7 = frontend_io_out_1_bits_cf_intrVec_7; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire  _T_6_T_29_cf_intrVec_8 = frontend_io_out_1_bits_cf_intrVec_8; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire  _T_6_T_29_cf_intrVec_9 = frontend_io_out_1_bits_cf_intrVec_9; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire  _T_6_T_29_cf_intrVec_10 = frontend_io_out_1_bits_cf_intrVec_10; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire  _T_6_T_29_cf_intrVec_11 = frontend_io_out_1_bits_cf_intrVec_11; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire [1:0] _T_31 = _T_7 + _T_19; // @[PipelineVector.scala 47:42]
  wire  _T_32 = ~frontend_io_out_0_valid; // @[PipelineVector.scala 50:39]
  wire [63:0] _GEN_1261 = 2'h1 == _T_8 ? _T_6_1_cf_instr : _T_6_0_cf_instr; // @[PipelineVector.scala 55:15]
  wire [38:0] _GEN_1262 = 2'h1 == _T_8 ? _T_6_1_cf_pc : _T_6_0_cf_pc; // @[PipelineVector.scala 55:15]
  wire [38:0] _GEN_1263 = 2'h1 == _T_8 ? _T_6_1_cf_pnpc : _T_6_0_cf_pnpc; // @[PipelineVector.scala 55:15]
  wire  _GEN_1268 = 2'h1 == _T_8 ? _T_6_1_cf_exceptionVec_1 : _T_6_0_cf_exceptionVec_1; // @[PipelineVector.scala 55:15]
  wire  _GEN_1269 = 2'h1 == _T_8 ? _T_6_1_cf_exceptionVec_2 : _T_6_0_cf_exceptionVec_2; // @[PipelineVector.scala 55:15]
  wire  _GEN_1279 = 2'h1 == _T_8 ? _T_6_1_cf_exceptionVec_12 : _T_6_0_cf_exceptionVec_12; // @[PipelineVector.scala 55:15]
  wire  _GEN_1283 = 2'h1 == _T_8 ? _T_6_1_cf_intrVec_0 : _T_6_0_cf_intrVec_0; // @[PipelineVector.scala 55:15]
  wire  _GEN_1284 = 2'h1 == _T_8 ? _T_6_1_cf_intrVec_1 : _T_6_0_cf_intrVec_1; // @[PipelineVector.scala 55:15]
  wire  _GEN_1285 = 2'h1 == _T_8 ? _T_6_1_cf_intrVec_2 : _T_6_0_cf_intrVec_2; // @[PipelineVector.scala 55:15]
  wire  _GEN_1286 = 2'h1 == _T_8 ? _T_6_1_cf_intrVec_3 : _T_6_0_cf_intrVec_3; // @[PipelineVector.scala 55:15]
  wire  _GEN_1287 = 2'h1 == _T_8 ? _T_6_1_cf_intrVec_4 : _T_6_0_cf_intrVec_4; // @[PipelineVector.scala 55:15]
  wire  _GEN_1288 = 2'h1 == _T_8 ? _T_6_1_cf_intrVec_5 : _T_6_0_cf_intrVec_5; // @[PipelineVector.scala 55:15]
  wire  _GEN_1289 = 2'h1 == _T_8 ? _T_6_1_cf_intrVec_6 : _T_6_0_cf_intrVec_6; // @[PipelineVector.scala 55:15]
  wire  _GEN_1290 = 2'h1 == _T_8 ? _T_6_1_cf_intrVec_7 : _T_6_0_cf_intrVec_7; // @[PipelineVector.scala 55:15]
  wire  _GEN_1291 = 2'h1 == _T_8 ? _T_6_1_cf_intrVec_8 : _T_6_0_cf_intrVec_8; // @[PipelineVector.scala 55:15]
  wire  _GEN_1292 = 2'h1 == _T_8 ? _T_6_1_cf_intrVec_9 : _T_6_0_cf_intrVec_9; // @[PipelineVector.scala 55:15]
  wire  _GEN_1293 = 2'h1 == _T_8 ? _T_6_1_cf_intrVec_10 : _T_6_0_cf_intrVec_10; // @[PipelineVector.scala 55:15]
  wire  _GEN_1294 = 2'h1 == _T_8 ? _T_6_1_cf_intrVec_11 : _T_6_0_cf_intrVec_11; // @[PipelineVector.scala 55:15]
  wire [3:0] _GEN_1295 = 2'h1 == _T_8 ? _T_6_1_cf_brIdx : _T_6_0_cf_brIdx; // @[PipelineVector.scala 55:15]
  wire  _GEN_1297 = 2'h1 == _T_8 ? _T_6_1_cf_crossPageIPFFix : _T_6_0_cf_crossPageIPFFix; // @[PipelineVector.scala 55:15]
  wire [1:0] _GEN_1298 = 2'h1 == _T_8 ? _T_6_1_ctrl_src1Type : _T_6_0_ctrl_src1Type; // @[PipelineVector.scala 55:15]
  wire [1:0] _GEN_1299 = 2'h1 == _T_8 ? _T_6_1_ctrl_src2Type : _T_6_0_ctrl_src2Type; // @[PipelineVector.scala 55:15]
  wire [2:0] _GEN_1300 = 2'h1 == _T_8 ? _T_6_1_ctrl_fuType : _T_6_0_ctrl_fuType; // @[PipelineVector.scala 55:15]
  wire [6:0] _GEN_1301 = 2'h1 == _T_8 ? _T_6_1_ctrl_fuOpType : _T_6_0_ctrl_fuOpType; // @[PipelineVector.scala 55:15]
  wire [4:0] _GEN_1302 = 2'h1 == _T_8 ? _T_6_1_ctrl_rfSrc1 : _T_6_0_ctrl_rfSrc1; // @[PipelineVector.scala 55:15]
  wire [4:0] _GEN_1303 = 2'h1 == _T_8 ? _T_6_1_ctrl_rfSrc2 : _T_6_0_ctrl_rfSrc2; // @[PipelineVector.scala 55:15]
  wire  _GEN_1304 = 2'h1 == _T_8 ? _T_6_1_ctrl_rfWen : _T_6_0_ctrl_rfWen; // @[PipelineVector.scala 55:15]
  wire [4:0] _GEN_1305 = 2'h1 == _T_8 ? _T_6_1_ctrl_rfDest : _T_6_0_ctrl_rfDest; // @[PipelineVector.scala 55:15]
  wire  _GEN_1308 = 2'h1 == _T_8 ? _T_6_1_ctrl_isNutCoreTrap : _T_6_0_ctrl_isNutCoreTrap; // @[PipelineVector.scala 55:15]
  wire [63:0] _GEN_1315 = 2'h1 == _T_8 ? _T_6_1_data_imm : _T_6_0_data_imm; // @[PipelineVector.scala 55:15]
  wire [63:0] _GEN_1321 = 2'h2 == _T_8 ? _T_6_2_cf_instr : _GEN_1261; // @[PipelineVector.scala 55:15]
  wire [38:0] _GEN_1322 = 2'h2 == _T_8 ? _T_6_2_cf_pc : _GEN_1262; // @[PipelineVector.scala 55:15]
  wire [38:0] _GEN_1323 = 2'h2 == _T_8 ? _T_6_2_cf_pnpc : _GEN_1263; // @[PipelineVector.scala 55:15]
  wire  _GEN_1328 = 2'h2 == _T_8 ? _T_6_2_cf_exceptionVec_1 : _GEN_1268; // @[PipelineVector.scala 55:15]
  wire  _GEN_1329 = 2'h2 == _T_8 ? _T_6_2_cf_exceptionVec_2 : _GEN_1269; // @[PipelineVector.scala 55:15]
  wire  _GEN_1339 = 2'h2 == _T_8 ? _T_6_2_cf_exceptionVec_12 : _GEN_1279; // @[PipelineVector.scala 55:15]
  wire  _GEN_1343 = 2'h2 == _T_8 ? _T_6_2_cf_intrVec_0 : _GEN_1283; // @[PipelineVector.scala 55:15]
  wire  _GEN_1344 = 2'h2 == _T_8 ? _T_6_2_cf_intrVec_1 : _GEN_1284; // @[PipelineVector.scala 55:15]
  wire  _GEN_1345 = 2'h2 == _T_8 ? _T_6_2_cf_intrVec_2 : _GEN_1285; // @[PipelineVector.scala 55:15]
  wire  _GEN_1346 = 2'h2 == _T_8 ? _T_6_2_cf_intrVec_3 : _GEN_1286; // @[PipelineVector.scala 55:15]
  wire  _GEN_1347 = 2'h2 == _T_8 ? _T_6_2_cf_intrVec_4 : _GEN_1287; // @[PipelineVector.scala 55:15]
  wire  _GEN_1348 = 2'h2 == _T_8 ? _T_6_2_cf_intrVec_5 : _GEN_1288; // @[PipelineVector.scala 55:15]
  wire  _GEN_1349 = 2'h2 == _T_8 ? _T_6_2_cf_intrVec_6 : _GEN_1289; // @[PipelineVector.scala 55:15]
  wire  _GEN_1350 = 2'h2 == _T_8 ? _T_6_2_cf_intrVec_7 : _GEN_1290; // @[PipelineVector.scala 55:15]
  wire  _GEN_1351 = 2'h2 == _T_8 ? _T_6_2_cf_intrVec_8 : _GEN_1291; // @[PipelineVector.scala 55:15]
  wire  _GEN_1352 = 2'h2 == _T_8 ? _T_6_2_cf_intrVec_9 : _GEN_1292; // @[PipelineVector.scala 55:15]
  wire  _GEN_1353 = 2'h2 == _T_8 ? _T_6_2_cf_intrVec_10 : _GEN_1293; // @[PipelineVector.scala 55:15]
  wire  _GEN_1354 = 2'h2 == _T_8 ? _T_6_2_cf_intrVec_11 : _GEN_1294; // @[PipelineVector.scala 55:15]
  wire [3:0] _GEN_1355 = 2'h2 == _T_8 ? _T_6_2_cf_brIdx : _GEN_1295; // @[PipelineVector.scala 55:15]
  wire  _GEN_1357 = 2'h2 == _T_8 ? _T_6_2_cf_crossPageIPFFix : _GEN_1297; // @[PipelineVector.scala 55:15]
  wire [1:0] _GEN_1358 = 2'h2 == _T_8 ? _T_6_2_ctrl_src1Type : _GEN_1298; // @[PipelineVector.scala 55:15]
  wire [1:0] _GEN_1359 = 2'h2 == _T_8 ? _T_6_2_ctrl_src2Type : _GEN_1299; // @[PipelineVector.scala 55:15]
  wire [2:0] _GEN_1360 = 2'h2 == _T_8 ? _T_6_2_ctrl_fuType : _GEN_1300; // @[PipelineVector.scala 55:15]
  wire [6:0] _GEN_1361 = 2'h2 == _T_8 ? _T_6_2_ctrl_fuOpType : _GEN_1301; // @[PipelineVector.scala 55:15]
  wire [4:0] _GEN_1362 = 2'h2 == _T_8 ? _T_6_2_ctrl_rfSrc1 : _GEN_1302; // @[PipelineVector.scala 55:15]
  wire [4:0] _GEN_1363 = 2'h2 == _T_8 ? _T_6_2_ctrl_rfSrc2 : _GEN_1303; // @[PipelineVector.scala 55:15]
  wire  _GEN_1364 = 2'h2 == _T_8 ? _T_6_2_ctrl_rfWen : _GEN_1304; // @[PipelineVector.scala 55:15]
  wire [4:0] _GEN_1365 = 2'h2 == _T_8 ? _T_6_2_ctrl_rfDest : _GEN_1305; // @[PipelineVector.scala 55:15]
  wire  _GEN_1368 = 2'h2 == _T_8 ? _T_6_2_ctrl_isNutCoreTrap : _GEN_1308; // @[PipelineVector.scala 55:15]
  wire [63:0] _GEN_1375 = 2'h2 == _T_8 ? _T_6_2_data_imm : _GEN_1315; // @[PipelineVector.scala 55:15]
  wire  _T_41 = Backend_inorder_io_in_0_ready & Backend_inorder_io_in_0_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _T_43 = {{1'd0}, _T_41}; // @[PipelineVector.scala 64:44]
  wire  _T_44 = _T_43 > 2'h0; // @[PipelineVector.scala 65:35]
  wire [1:0] _T_46 = _T_8 + _T_43; // @[PipelineVector.scala 67:42]
  wire [3:0] _T_49 = 3'h4 + _T_25; // @[PipelineVector.scala 77:86]
  wire [3:0] _GEN_1685 = {{2'd0}, _T_8}; // @[PipelineVector.scala 77:113]
  wire [3:0] _T_51 = _T_49 - _GEN_1685; // @[PipelineVector.scala 77:113]
  wire [3:0] _GEN_0 = _T_51 % 4'h4; // @[PipelineVector.scala 77:140]
  wire [2:0] _T_52 = _GEN_0[2:0]; // @[PipelineVector.scala 77:140]
  wire  _T_54 = ~reset; // @[PipelineVector.scala 77:15]
  reg [63:0] _T_62; // @[GTimer.scala 24:20]
  wire [63:0] _T_64 = _T_62 + 64'h1; // @[GTimer.scala 25:12]
  Frontend_inorder frontend ( // @[NutCore.scala 102:34]
    .clock(frontend_clock),
    .reset(frontend_reset),
    .io_out_0_ready(frontend_io_out_0_ready),
    .io_out_0_valid(frontend_io_out_0_valid),
    .io_out_0_bits_cf_instr(frontend_io_out_0_bits_cf_instr),
    .io_out_0_bits_cf_pc(frontend_io_out_0_bits_cf_pc),
    .io_out_0_bits_cf_pnpc(frontend_io_out_0_bits_cf_pnpc),
    .io_out_0_bits_cf_exceptionVec_1(frontend_io_out_0_bits_cf_exceptionVec_1),
    .io_out_0_bits_cf_exceptionVec_2(frontend_io_out_0_bits_cf_exceptionVec_2),
    .io_out_0_bits_cf_exceptionVec_12(frontend_io_out_0_bits_cf_exceptionVec_12),
    .io_out_0_bits_cf_intrVec_0(frontend_io_out_0_bits_cf_intrVec_0),
    .io_out_0_bits_cf_intrVec_1(frontend_io_out_0_bits_cf_intrVec_1),
    .io_out_0_bits_cf_intrVec_2(frontend_io_out_0_bits_cf_intrVec_2),
    .io_out_0_bits_cf_intrVec_3(frontend_io_out_0_bits_cf_intrVec_3),
    .io_out_0_bits_cf_intrVec_4(frontend_io_out_0_bits_cf_intrVec_4),
    .io_out_0_bits_cf_intrVec_5(frontend_io_out_0_bits_cf_intrVec_5),
    .io_out_0_bits_cf_intrVec_6(frontend_io_out_0_bits_cf_intrVec_6),
    .io_out_0_bits_cf_intrVec_7(frontend_io_out_0_bits_cf_intrVec_7),
    .io_out_0_bits_cf_intrVec_8(frontend_io_out_0_bits_cf_intrVec_8),
    .io_out_0_bits_cf_intrVec_9(frontend_io_out_0_bits_cf_intrVec_9),
    .io_out_0_bits_cf_intrVec_10(frontend_io_out_0_bits_cf_intrVec_10),
    .io_out_0_bits_cf_intrVec_11(frontend_io_out_0_bits_cf_intrVec_11),
    .io_out_0_bits_cf_brIdx(frontend_io_out_0_bits_cf_brIdx),
    .io_out_0_bits_cf_crossPageIPFFix(frontend_io_out_0_bits_cf_crossPageIPFFix),
    .io_out_0_bits_ctrl_src1Type(frontend_io_out_0_bits_ctrl_src1Type),
    .io_out_0_bits_ctrl_src2Type(frontend_io_out_0_bits_ctrl_src2Type),
    .io_out_0_bits_ctrl_fuType(frontend_io_out_0_bits_ctrl_fuType),
    .io_out_0_bits_ctrl_fuOpType(frontend_io_out_0_bits_ctrl_fuOpType),
    .io_out_0_bits_ctrl_rfSrc1(frontend_io_out_0_bits_ctrl_rfSrc1),
    .io_out_0_bits_ctrl_rfSrc2(frontend_io_out_0_bits_ctrl_rfSrc2),
    .io_out_0_bits_ctrl_rfWen(frontend_io_out_0_bits_ctrl_rfWen),
    .io_out_0_bits_ctrl_rfDest(frontend_io_out_0_bits_ctrl_rfDest),
    .io_out_0_bits_ctrl_isNutCoreTrap(frontend_io_out_0_bits_ctrl_isNutCoreTrap),
    .io_out_0_bits_data_imm(frontend_io_out_0_bits_data_imm),
    .io_out_1_bits_cf_intrVec_0(frontend_io_out_1_bits_cf_intrVec_0),
    .io_out_1_bits_cf_intrVec_1(frontend_io_out_1_bits_cf_intrVec_1),
    .io_out_1_bits_cf_intrVec_2(frontend_io_out_1_bits_cf_intrVec_2),
    .io_out_1_bits_cf_intrVec_3(frontend_io_out_1_bits_cf_intrVec_3),
    .io_out_1_bits_cf_intrVec_4(frontend_io_out_1_bits_cf_intrVec_4),
    .io_out_1_bits_cf_intrVec_5(frontend_io_out_1_bits_cf_intrVec_5),
    .io_out_1_bits_cf_intrVec_6(frontend_io_out_1_bits_cf_intrVec_6),
    .io_out_1_bits_cf_intrVec_7(frontend_io_out_1_bits_cf_intrVec_7),
    .io_out_1_bits_cf_intrVec_8(frontend_io_out_1_bits_cf_intrVec_8),
    .io_out_1_bits_cf_intrVec_9(frontend_io_out_1_bits_cf_intrVec_9),
    .io_out_1_bits_cf_intrVec_10(frontend_io_out_1_bits_cf_intrVec_10),
    .io_out_1_bits_cf_intrVec_11(frontend_io_out_1_bits_cf_intrVec_11),
    .io_imem_req_ready(frontend_io_imem_req_ready),
    .io_imem_req_valid(frontend_io_imem_req_valid),
    .io_imem_req_bits_addr(frontend_io_imem_req_bits_addr),
    .io_imem_req_bits_user(frontend_io_imem_req_bits_user),
    .io_imem_resp_ready(frontend_io_imem_resp_ready),
    .io_imem_resp_valid(frontend_io_imem_resp_valid),
    .io_imem_resp_bits_rdata(frontend_io_imem_resp_bits_rdata),
    .io_imem_resp_bits_user(frontend_io_imem_resp_bits_user),
    .io_flushVec(frontend_io_flushVec),
    .io_ipf(frontend_io_ipf),
    .io_redirect_target(frontend_io_redirect_target),
    .io_redirect_valid(frontend_io_redirect_valid),
    .flushICache(frontend_flushICache),
    ._T_243_valid(frontend__T_243_valid),
    ._T_243_pc(frontend__T_243_pc),
    ._T_243_isMissPredict(frontend__T_243_isMissPredict),
    ._T_243_actualTarget(frontend__T_243_actualTarget),
    ._T_243_actualTaken(frontend__T_243_actualTaken),
    ._T_243_fuOpType(frontend__T_243_fuOpType),
    ._T_243_btbType(frontend__T_243_btbType),
    ._T_243_isRVC(frontend__T_243_isRVC),
    .DISPLAY_ENABLE(frontend_DISPLAY_ENABLE),
    .vmEnable(frontend_vmEnable),
    .intrVec(frontend_intrVec),
    ._T_0(frontend__T_0),
    ._T_65(frontend__T_65),
    .flushTLB(frontend_flushTLB),
    ._T_66(frontend__T_66)
  );
  Backend_inorder Backend_inorder ( // @[NutCore.scala 144:25]
    .clock(Backend_inorder_clock),
    .reset(Backend_inorder_reset),
    .io_in_0_ready(Backend_inorder_io_in_0_ready),
    .io_in_0_valid(Backend_inorder_io_in_0_valid),
    .io_in_0_bits_cf_instr(Backend_inorder_io_in_0_bits_cf_instr),
    .io_in_0_bits_cf_pc(Backend_inorder_io_in_0_bits_cf_pc),
    .io_in_0_bits_cf_pnpc(Backend_inorder_io_in_0_bits_cf_pnpc),
    .io_in_0_bits_cf_exceptionVec_1(Backend_inorder_io_in_0_bits_cf_exceptionVec_1),
    .io_in_0_bits_cf_exceptionVec_2(Backend_inorder_io_in_0_bits_cf_exceptionVec_2),
    .io_in_0_bits_cf_exceptionVec_12(Backend_inorder_io_in_0_bits_cf_exceptionVec_12),
    .io_in_0_bits_cf_intrVec_0(Backend_inorder_io_in_0_bits_cf_intrVec_0),
    .io_in_0_bits_cf_intrVec_1(Backend_inorder_io_in_0_bits_cf_intrVec_1),
    .io_in_0_bits_cf_intrVec_2(Backend_inorder_io_in_0_bits_cf_intrVec_2),
    .io_in_0_bits_cf_intrVec_3(Backend_inorder_io_in_0_bits_cf_intrVec_3),
    .io_in_0_bits_cf_intrVec_4(Backend_inorder_io_in_0_bits_cf_intrVec_4),
    .io_in_0_bits_cf_intrVec_5(Backend_inorder_io_in_0_bits_cf_intrVec_5),
    .io_in_0_bits_cf_intrVec_6(Backend_inorder_io_in_0_bits_cf_intrVec_6),
    .io_in_0_bits_cf_intrVec_7(Backend_inorder_io_in_0_bits_cf_intrVec_7),
    .io_in_0_bits_cf_intrVec_8(Backend_inorder_io_in_0_bits_cf_intrVec_8),
    .io_in_0_bits_cf_intrVec_9(Backend_inorder_io_in_0_bits_cf_intrVec_9),
    .io_in_0_bits_cf_intrVec_10(Backend_inorder_io_in_0_bits_cf_intrVec_10),
    .io_in_0_bits_cf_intrVec_11(Backend_inorder_io_in_0_bits_cf_intrVec_11),
    .io_in_0_bits_cf_brIdx(Backend_inorder_io_in_0_bits_cf_brIdx),
    .io_in_0_bits_cf_crossPageIPFFix(Backend_inorder_io_in_0_bits_cf_crossPageIPFFix),
    .io_in_0_bits_ctrl_src1Type(Backend_inorder_io_in_0_bits_ctrl_src1Type),
    .io_in_0_bits_ctrl_src2Type(Backend_inorder_io_in_0_bits_ctrl_src2Type),
    .io_in_0_bits_ctrl_fuType(Backend_inorder_io_in_0_bits_ctrl_fuType),
    .io_in_0_bits_ctrl_fuOpType(Backend_inorder_io_in_0_bits_ctrl_fuOpType),
    .io_in_0_bits_ctrl_rfSrc1(Backend_inorder_io_in_0_bits_ctrl_rfSrc1),
    .io_in_0_bits_ctrl_rfSrc2(Backend_inorder_io_in_0_bits_ctrl_rfSrc2),
    .io_in_0_bits_ctrl_rfWen(Backend_inorder_io_in_0_bits_ctrl_rfWen),
    .io_in_0_bits_ctrl_rfDest(Backend_inorder_io_in_0_bits_ctrl_rfDest),
    .io_in_0_bits_ctrl_isNutCoreTrap(Backend_inorder_io_in_0_bits_ctrl_isNutCoreTrap),
    .io_in_0_bits_data_imm(Backend_inorder_io_in_0_bits_data_imm),
    .io_flush(Backend_inorder_io_flush),
    .io_dmem_req_ready(Backend_inorder_io_dmem_req_ready),
    .io_dmem_req_valid(Backend_inorder_io_dmem_req_valid),
    .io_dmem_req_bits_addr(Backend_inorder_io_dmem_req_bits_addr),
    .io_dmem_req_bits_size(Backend_inorder_io_dmem_req_bits_size),
    .io_dmem_req_bits_cmd(Backend_inorder_io_dmem_req_bits_cmd),
    .io_dmem_req_bits_wmask(Backend_inorder_io_dmem_req_bits_wmask),
    .io_dmem_req_bits_wdata(Backend_inorder_io_dmem_req_bits_wdata),
    .io_dmem_resp_valid(Backend_inorder_io_dmem_resp_valid),
    .io_dmem_resp_bits_rdata(Backend_inorder_io_dmem_resp_bits_rdata),
    .io_memMMU_imem_priviledgeMode(Backend_inorder_io_memMMU_imem_priviledgeMode),
    .io_memMMU_dmem_priviledgeMode(Backend_inorder_io_memMMU_dmem_priviledgeMode),
    .io_memMMU_dmem_status_sum(Backend_inorder_io_memMMU_dmem_status_sum),
    .io_memMMU_dmem_status_mxr(Backend_inorder_io_memMMU_dmem_status_mxr),
    .io_memMMU_dmem_loadPF(Backend_inorder_io_memMMU_dmem_loadPF),
    .io_memMMU_dmem_storePF(Backend_inorder_io_memMMU_dmem_storePF),
    .io_memMMU_dmem_addr(Backend_inorder_io_memMMU_dmem_addr),
    .io_redirect_target(Backend_inorder_io_redirect_target),
    .io_redirect_valid(Backend_inorder_io_redirect_valid),
    ._T_4181(Backend_inorder__T_4181),
    ._T_4184(Backend_inorder__T_4184),
    ._T_38(Backend_inorder__T_38),
    .flushICache(Backend_inorder_flushICache),
    ._T_4185(Backend_inorder__T_4185),
    .falseWire(Backend_inorder_falseWire),
    .satp(Backend_inorder_satp),
    ._T_243_valid(Backend_inorder__T_243_valid),
    ._T_243_pc(Backend_inorder__T_243_pc),
    ._T_243_isMissPredict(Backend_inorder__T_243_isMissPredict),
    ._T_243_actualTarget(Backend_inorder__T_243_actualTarget),
    ._T_243_actualTaken(Backend_inorder__T_243_actualTaken),
    ._T_243_fuOpType(Backend_inorder__T_243_fuOpType),
    ._T_243_btbType(Backend_inorder__T_243_btbType),
    ._T_243_isRVC(Backend_inorder__T_243_isRVC),
    .falseWire_0(Backend_inorder_falseWire_0),
    ._T_4178(Backend_inorder__T_4178),
    ._T_284_0(Backend_inorder__T_284_0),
    ._T_284_1(Backend_inorder__T_284_1),
    ._T_284_2(Backend_inorder__T_284_2),
    ._T_284_3(Backend_inorder__T_284_3),
    ._T_284_4(Backend_inorder__T_284_4),
    ._T_284_5(Backend_inorder__T_284_5),
    ._T_284_6(Backend_inorder__T_284_6),
    ._T_284_7(Backend_inorder__T_284_7),
    ._T_284_8(Backend_inorder__T_284_8),
    ._T_284_9(Backend_inorder__T_284_9),
    ._T_284_10(Backend_inorder__T_284_10),
    ._T_284_11(Backend_inorder__T_284_11),
    ._T_284_12(Backend_inorder__T_284_12),
    ._T_284_13(Backend_inorder__T_284_13),
    ._T_284_14(Backend_inorder__T_284_14),
    ._T_284_15(Backend_inorder__T_284_15),
    ._T_284_16(Backend_inorder__T_284_16),
    ._T_284_17(Backend_inorder__T_284_17),
    ._T_284_18(Backend_inorder__T_284_18),
    ._T_284_19(Backend_inorder__T_284_19),
    ._T_284_20(Backend_inorder__T_284_20),
    ._T_284_21(Backend_inorder__T_284_21),
    ._T_284_22(Backend_inorder__T_284_22),
    ._T_284_23(Backend_inorder__T_284_23),
    ._T_284_24(Backend_inorder__T_284_24),
    ._T_284_25(Backend_inorder__T_284_25),
    ._T_284_26(Backend_inorder__T_284_26),
    ._T_284_27(Backend_inorder__T_284_27),
    ._T_284_28(Backend_inorder__T_284_28),
    ._T_284_29(Backend_inorder__T_284_29),
    ._T_284_30(Backend_inorder__T_284_30),
    ._T_284_31(Backend_inorder__T_284_31),
    .mmio(Backend_inorder_mmio),
    ._T_36(Backend_inorder__T_36),
    .io_extra_mtip(Backend_inorder_io_extra_mtip),
    .amoReq(Backend_inorder_amoReq),
    ._T_32(Backend_inorder__T_32),
    ._T_13(Backend_inorder__T_13),
    .io_extra_meip_0(Backend_inorder_io_extra_meip_0),
    .vmEnable(Backend_inorder_vmEnable),
    ._T_31(Backend_inorder__T_31),
    ._T_37(Backend_inorder__T_37),
    ._T_26(Backend_inorder__T_26),
    .intrVec(Backend_inorder_intrVec),
    ._T_37_0(Backend_inorder__T_37_0),
    .io_extra_msip(Backend_inorder_io_extra_msip),
    ._T_65(Backend_inorder__T_65),
    ._T_4183(Backend_inorder__T_4183),
    ._T_4182(Backend_inorder__T_4182),
    .flushTLB(Backend_inorder_flushTLB),
    ._T_33(Backend_inorder__T_33),
    ._T_66(Backend_inorder__T_66),
    ._T_4179(Backend_inorder__T_4179)
  );
  SimpleBusCrossbarNto1 SimpleBusCrossbarNto1 ( // @[NutCore.scala 148:26]
    .clock(SimpleBusCrossbarNto1_clock),
    .reset(SimpleBusCrossbarNto1_reset),
    .io_in_0_req_ready(SimpleBusCrossbarNto1_io_in_0_req_ready),
    .io_in_0_req_valid(SimpleBusCrossbarNto1_io_in_0_req_valid),
    .io_in_0_req_bits_addr(SimpleBusCrossbarNto1_io_in_0_req_bits_addr),
    .io_in_0_req_bits_cmd(SimpleBusCrossbarNto1_io_in_0_req_bits_cmd),
    .io_in_0_req_bits_wmask(SimpleBusCrossbarNto1_io_in_0_req_bits_wmask),
    .io_in_0_req_bits_wdata(SimpleBusCrossbarNto1_io_in_0_req_bits_wdata),
    .io_in_0_resp_valid(SimpleBusCrossbarNto1_io_in_0_resp_valid),
    .io_in_0_resp_bits_cmd(SimpleBusCrossbarNto1_io_in_0_resp_bits_cmd),
    .io_in_0_resp_bits_rdata(SimpleBusCrossbarNto1_io_in_0_resp_bits_rdata),
    .io_in_1_req_ready(SimpleBusCrossbarNto1_io_in_1_req_ready),
    .io_in_1_req_valid(SimpleBusCrossbarNto1_io_in_1_req_valid),
    .io_in_1_req_bits_addr(SimpleBusCrossbarNto1_io_in_1_req_bits_addr),
    .io_in_1_req_bits_size(SimpleBusCrossbarNto1_io_in_1_req_bits_size),
    .io_in_1_req_bits_cmd(SimpleBusCrossbarNto1_io_in_1_req_bits_cmd),
    .io_in_1_req_bits_wmask(SimpleBusCrossbarNto1_io_in_1_req_bits_wmask),
    .io_in_1_req_bits_wdata(SimpleBusCrossbarNto1_io_in_1_req_bits_wdata),
    .io_in_1_resp_valid(SimpleBusCrossbarNto1_io_in_1_resp_valid),
    .io_in_1_resp_bits_cmd(SimpleBusCrossbarNto1_io_in_1_resp_bits_cmd),
    .io_in_1_resp_bits_rdata(SimpleBusCrossbarNto1_io_in_1_resp_bits_rdata),
    .io_out_req_ready(SimpleBusCrossbarNto1_io_out_req_ready),
    .io_out_req_valid(SimpleBusCrossbarNto1_io_out_req_valid),
    .io_out_req_bits_addr(SimpleBusCrossbarNto1_io_out_req_bits_addr),
    .io_out_req_bits_size(SimpleBusCrossbarNto1_io_out_req_bits_size),
    .io_out_req_bits_cmd(SimpleBusCrossbarNto1_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(SimpleBusCrossbarNto1_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(SimpleBusCrossbarNto1_io_out_req_bits_wdata),
    .io_out_resp_ready(SimpleBusCrossbarNto1_io_out_resp_ready),
    .io_out_resp_valid(SimpleBusCrossbarNto1_io_out_resp_valid),
    .io_out_resp_bits_cmd(SimpleBusCrossbarNto1_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(SimpleBusCrossbarNto1_io_out_resp_bits_rdata)
  );
  SimpleBusCrossbarNto1_1 SimpleBusCrossbarNto1_1 ( // @[NutCore.scala 149:26]
    .clock(SimpleBusCrossbarNto1_1_clock),
    .reset(SimpleBusCrossbarNto1_1_reset),
    .io_in_0_req_ready(SimpleBusCrossbarNto1_1_io_in_0_req_ready),
    .io_in_0_req_valid(SimpleBusCrossbarNto1_1_io_in_0_req_valid),
    .io_in_0_req_bits_addr(SimpleBusCrossbarNto1_1_io_in_0_req_bits_addr),
    .io_in_0_req_bits_size(SimpleBusCrossbarNto1_1_io_in_0_req_bits_size),
    .io_in_0_req_bits_cmd(SimpleBusCrossbarNto1_1_io_in_0_req_bits_cmd),
    .io_in_0_req_bits_wmask(SimpleBusCrossbarNto1_1_io_in_0_req_bits_wmask),
    .io_in_0_req_bits_wdata(SimpleBusCrossbarNto1_1_io_in_0_req_bits_wdata),
    .io_in_0_resp_valid(SimpleBusCrossbarNto1_1_io_in_0_resp_valid),
    .io_in_0_resp_bits_cmd(SimpleBusCrossbarNto1_1_io_in_0_resp_bits_cmd),
    .io_in_0_resp_bits_rdata(SimpleBusCrossbarNto1_1_io_in_0_resp_bits_rdata),
    .io_in_1_req_ready(SimpleBusCrossbarNto1_1_io_in_1_req_ready),
    .io_in_1_req_valid(SimpleBusCrossbarNto1_1_io_in_1_req_valid),
    .io_in_1_req_bits_addr(SimpleBusCrossbarNto1_1_io_in_1_req_bits_addr),
    .io_in_1_req_bits_cmd(SimpleBusCrossbarNto1_1_io_in_1_req_bits_cmd),
    .io_in_1_req_bits_wdata(SimpleBusCrossbarNto1_1_io_in_1_req_bits_wdata),
    .io_in_1_resp_valid(SimpleBusCrossbarNto1_1_io_in_1_resp_valid),
    .io_in_1_resp_bits_cmd(SimpleBusCrossbarNto1_1_io_in_1_resp_bits_cmd),
    .io_in_1_resp_bits_rdata(SimpleBusCrossbarNto1_1_io_in_1_resp_bits_rdata),
    .io_in_2_req_ready(SimpleBusCrossbarNto1_1_io_in_2_req_ready),
    .io_in_2_req_valid(SimpleBusCrossbarNto1_1_io_in_2_req_valid),
    .io_in_2_req_bits_addr(SimpleBusCrossbarNto1_1_io_in_2_req_bits_addr),
    .io_in_2_req_bits_cmd(SimpleBusCrossbarNto1_1_io_in_2_req_bits_cmd),
    .io_in_2_req_bits_wdata(SimpleBusCrossbarNto1_1_io_in_2_req_bits_wdata),
    .io_in_2_resp_valid(SimpleBusCrossbarNto1_1_io_in_2_resp_valid),
    .io_in_2_resp_bits_cmd(SimpleBusCrossbarNto1_1_io_in_2_resp_bits_cmd),
    .io_in_2_resp_bits_rdata(SimpleBusCrossbarNto1_1_io_in_2_resp_bits_rdata),
    .io_in_3_req_ready(SimpleBusCrossbarNto1_1_io_in_3_req_ready),
    .io_in_3_req_valid(SimpleBusCrossbarNto1_1_io_in_3_req_valid),
    .io_in_3_req_bits_addr(SimpleBusCrossbarNto1_1_io_in_3_req_bits_addr),
    .io_in_3_req_bits_size(SimpleBusCrossbarNto1_1_io_in_3_req_bits_size),
    .io_in_3_req_bits_cmd(SimpleBusCrossbarNto1_1_io_in_3_req_bits_cmd),
    .io_in_3_req_bits_wmask(SimpleBusCrossbarNto1_1_io_in_3_req_bits_wmask),
    .io_in_3_req_bits_wdata(SimpleBusCrossbarNto1_1_io_in_3_req_bits_wdata),
    .io_in_3_resp_ready(SimpleBusCrossbarNto1_1_io_in_3_resp_ready),
    .io_in_3_resp_valid(SimpleBusCrossbarNto1_1_io_in_3_resp_valid),
    .io_in_3_resp_bits_cmd(SimpleBusCrossbarNto1_1_io_in_3_resp_bits_cmd),
    .io_in_3_resp_bits_rdata(SimpleBusCrossbarNto1_1_io_in_3_resp_bits_rdata),
    .io_out_req_ready(SimpleBusCrossbarNto1_1_io_out_req_ready),
    .io_out_req_valid(SimpleBusCrossbarNto1_1_io_out_req_valid),
    .io_out_req_bits_addr(SimpleBusCrossbarNto1_1_io_out_req_bits_addr),
    .io_out_req_bits_size(SimpleBusCrossbarNto1_1_io_out_req_bits_size),
    .io_out_req_bits_cmd(SimpleBusCrossbarNto1_1_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(SimpleBusCrossbarNto1_1_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(SimpleBusCrossbarNto1_1_io_out_req_bits_wdata),
    .io_out_resp_ready(SimpleBusCrossbarNto1_1_io_out_resp_ready),
    .io_out_resp_valid(SimpleBusCrossbarNto1_1_io_out_resp_valid),
    .io_out_resp_bits_cmd(SimpleBusCrossbarNto1_1_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(SimpleBusCrossbarNto1_1_io_out_resp_bits_rdata)
  );
  EmbeddedTLB EmbeddedTLB ( // @[EmbeddedTLB.scala 427:23]
    .clock(EmbeddedTLB_clock),
    .reset(EmbeddedTLB_reset),
    .io_in_req_ready(EmbeddedTLB_io_in_req_ready),
    .io_in_req_valid(EmbeddedTLB_io_in_req_valid),
    .io_in_req_bits_addr(EmbeddedTLB_io_in_req_bits_addr),
    .io_in_req_bits_user(EmbeddedTLB_io_in_req_bits_user),
    .io_in_resp_ready(EmbeddedTLB_io_in_resp_ready),
    .io_in_resp_valid(EmbeddedTLB_io_in_resp_valid),
    .io_in_resp_bits_cmd(EmbeddedTLB_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(EmbeddedTLB_io_in_resp_bits_rdata),
    .io_in_resp_bits_user(EmbeddedTLB_io_in_resp_bits_user),
    .io_out_req_ready(EmbeddedTLB_io_out_req_ready),
    .io_out_req_valid(EmbeddedTLB_io_out_req_valid),
    .io_out_req_bits_addr(EmbeddedTLB_io_out_req_bits_addr),
    .io_out_req_bits_cmd(EmbeddedTLB_io_out_req_bits_cmd),
    .io_out_req_bits_wdata(EmbeddedTLB_io_out_req_bits_wdata),
    .io_out_req_bits_user(EmbeddedTLB_io_out_req_bits_user),
    .io_out_resp_ready(EmbeddedTLB_io_out_resp_ready),
    .io_out_resp_valid(EmbeddedTLB_io_out_resp_valid),
    .io_out_resp_bits_rdata(EmbeddedTLB_io_out_resp_bits_rdata),
    .io_out_resp_bits_user(EmbeddedTLB_io_out_resp_bits_user),
    .io_mem_req_ready(EmbeddedTLB_io_mem_req_ready),
    .io_mem_req_valid(EmbeddedTLB_io_mem_req_valid),
    .io_mem_req_bits_addr(EmbeddedTLB_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(EmbeddedTLB_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(EmbeddedTLB_io_mem_req_bits_wdata),
    .io_mem_resp_valid(EmbeddedTLB_io_mem_resp_valid),
    .io_mem_resp_bits_cmd(EmbeddedTLB_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_rdata(EmbeddedTLB_io_mem_resp_bits_rdata),
    .io_flush(EmbeddedTLB_io_flush),
    .io_csrMMU_priviledgeMode(EmbeddedTLB_io_csrMMU_priviledgeMode),
    .io_csrMMU_loadPF(EmbeddedTLB_io_csrMMU_loadPF),
    .io_csrMMU_storePF(EmbeddedTLB_io_csrMMU_storePF),
    .io_cacheEmpty(EmbeddedTLB_io_cacheEmpty),
    .io_ipf(EmbeddedTLB_io_ipf),
    .CSRSATP(EmbeddedTLB_CSRSATP),
    .DISPLAY_ENABLE(EmbeddedTLB_DISPLAY_ENABLE),
    .MOUFlushTLB(EmbeddedTLB_MOUFlushTLB)
  );
  Cache Cache ( // @[Cache.scala 678:35]
    .clock(Cache_clock),
    .reset(Cache_reset),
    .io_in_req_ready(Cache_io_in_req_ready),
    .io_in_req_valid(Cache_io_in_req_valid),
    .io_in_req_bits_addr(Cache_io_in_req_bits_addr),
    .io_in_req_bits_user(Cache_io_in_req_bits_user),
    .io_in_resp_ready(Cache_io_in_resp_ready),
    .io_in_resp_valid(Cache_io_in_resp_valid),
    .io_in_resp_bits_rdata(Cache_io_in_resp_bits_rdata),
    .io_in_resp_bits_user(Cache_io_in_resp_bits_user),
    .io_flush(Cache_io_flush),
    .io_out_mem_req_ready(Cache_io_out_mem_req_ready),
    .io_out_mem_req_valid(Cache_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(Cache_io_out_mem_req_bits_addr),
    .io_out_mem_req_bits_cmd(Cache_io_out_mem_req_bits_cmd),
    .io_out_mem_req_bits_wdata(Cache_io_out_mem_req_bits_wdata),
    .io_out_mem_resp_valid(Cache_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_cmd(Cache_io_out_mem_resp_bits_cmd),
    .io_out_mem_resp_bits_rdata(Cache_io_out_mem_resp_bits_rdata),
    .io_mmio_req_ready(Cache_io_mmio_req_ready),
    .io_mmio_req_valid(Cache_io_mmio_req_valid),
    .io_mmio_req_bits_addr(Cache_io_mmio_req_bits_addr),
    .io_mmio_resp_valid(Cache_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(Cache_io_mmio_resp_bits_rdata),
    .io_empty(Cache_io_empty),
    .MOUFlushICache(Cache_MOUFlushICache),
    .DISPLAY_ENABLE(Cache_DISPLAY_ENABLE)
  );
  EmbeddedTLB_1 EmbeddedTLB_1 ( // @[EmbeddedTLB.scala 427:23]
    .clock(EmbeddedTLB_1_clock),
    .reset(EmbeddedTLB_1_reset),
    .io_in_req_ready(EmbeddedTLB_1_io_in_req_ready),
    .io_in_req_valid(EmbeddedTLB_1_io_in_req_valid),
    .io_in_req_bits_addr(EmbeddedTLB_1_io_in_req_bits_addr),
    .io_in_req_bits_size(EmbeddedTLB_1_io_in_req_bits_size),
    .io_in_req_bits_cmd(EmbeddedTLB_1_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(EmbeddedTLB_1_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(EmbeddedTLB_1_io_in_req_bits_wdata),
    .io_in_resp_valid(EmbeddedTLB_1_io_in_resp_valid),
    .io_in_resp_bits_cmd(EmbeddedTLB_1_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(EmbeddedTLB_1_io_in_resp_bits_rdata),
    .io_out_req_ready(EmbeddedTLB_1_io_out_req_ready),
    .io_out_req_valid(EmbeddedTLB_1_io_out_req_valid),
    .io_out_req_bits_addr(EmbeddedTLB_1_io_out_req_bits_addr),
    .io_out_req_bits_size(EmbeddedTLB_1_io_out_req_bits_size),
    .io_out_req_bits_cmd(EmbeddedTLB_1_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(EmbeddedTLB_1_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(EmbeddedTLB_1_io_out_req_bits_wdata),
    .io_out_resp_ready(EmbeddedTLB_1_io_out_resp_ready),
    .io_out_resp_valid(EmbeddedTLB_1_io_out_resp_valid),
    .io_out_resp_bits_cmd(EmbeddedTLB_1_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(EmbeddedTLB_1_io_out_resp_bits_rdata),
    .io_mem_req_ready(EmbeddedTLB_1_io_mem_req_ready),
    .io_mem_req_valid(EmbeddedTLB_1_io_mem_req_valid),
    .io_mem_req_bits_addr(EmbeddedTLB_1_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(EmbeddedTLB_1_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(EmbeddedTLB_1_io_mem_req_bits_wdata),
    .io_mem_resp_valid(EmbeddedTLB_1_io_mem_resp_valid),
    .io_mem_resp_bits_cmd(EmbeddedTLB_1_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_rdata(EmbeddedTLB_1_io_mem_resp_bits_rdata),
    .io_csrMMU_priviledgeMode(EmbeddedTLB_1_io_csrMMU_priviledgeMode),
    .io_csrMMU_status_sum(EmbeddedTLB_1_io_csrMMU_status_sum),
    .io_csrMMU_status_mxr(EmbeddedTLB_1_io_csrMMU_status_mxr),
    .io_csrMMU_loadPF(EmbeddedTLB_1_io_csrMMU_loadPF),
    .io_csrMMU_storePF(EmbeddedTLB_1_io_csrMMU_storePF),
    .io_csrMMU_addr(EmbeddedTLB_1_io_csrMMU_addr),
    .io_cacheEmpty(EmbeddedTLB_1_io_cacheEmpty),
    .io_ipf(EmbeddedTLB_1_io_ipf),
    ._T_38_0(EmbeddedTLB_1__T_38_0),
    .CSRSATP(EmbeddedTLB_1_CSRSATP),
    .amoReq(EmbeddedTLB_1_amoReq),
    .DISPLAY_ENABLE(EmbeddedTLB_1_DISPLAY_ENABLE),
    .vmEnable_0(EmbeddedTLB_1_vmEnable_0),
    ._T_37_1(EmbeddedTLB_1__T_37_1),
    .MOUFlushTLB(EmbeddedTLB_1_MOUFlushTLB)
  );
  Cache_1 Cache_1 ( // @[Cache.scala 678:35]
    .clock(Cache_1_clock),
    .reset(Cache_1_reset),
    .io_in_req_ready(Cache_1_io_in_req_ready),
    .io_in_req_valid(Cache_1_io_in_req_valid),
    .io_in_req_bits_addr(Cache_1_io_in_req_bits_addr),
    .io_in_req_bits_size(Cache_1_io_in_req_bits_size),
    .io_in_req_bits_cmd(Cache_1_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(Cache_1_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(Cache_1_io_in_req_bits_wdata),
    .io_in_resp_ready(Cache_1_io_in_resp_ready),
    .io_in_resp_valid(Cache_1_io_in_resp_valid),
    .io_in_resp_bits_cmd(Cache_1_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(Cache_1_io_in_resp_bits_rdata),
    .io_out_mem_req_ready(Cache_1_io_out_mem_req_ready),
    .io_out_mem_req_valid(Cache_1_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(Cache_1_io_out_mem_req_bits_addr),
    .io_out_mem_req_bits_cmd(Cache_1_io_out_mem_req_bits_cmd),
    .io_out_mem_req_bits_wdata(Cache_1_io_out_mem_req_bits_wdata),
    .io_out_mem_resp_valid(Cache_1_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_cmd(Cache_1_io_out_mem_resp_bits_cmd),
    .io_out_mem_resp_bits_rdata(Cache_1_io_out_mem_resp_bits_rdata),
    .io_out_coh_req_ready(Cache_1_io_out_coh_req_ready),
    .io_out_coh_req_valid(Cache_1_io_out_coh_req_valid),
    .io_out_coh_req_bits_addr(Cache_1_io_out_coh_req_bits_addr),
    .io_out_coh_req_bits_wdata(Cache_1_io_out_coh_req_bits_wdata),
    .io_out_coh_resp_valid(Cache_1_io_out_coh_resp_valid),
    .io_out_coh_resp_bits_cmd(Cache_1_io_out_coh_resp_bits_cmd),
    .io_out_coh_resp_bits_rdata(Cache_1_io_out_coh_resp_bits_rdata),
    .io_mmio_req_ready(Cache_1_io_mmio_req_ready),
    .io_mmio_req_valid(Cache_1_io_mmio_req_valid),
    .io_mmio_req_bits_addr(Cache_1_io_mmio_req_bits_addr),
    .io_mmio_req_bits_size(Cache_1_io_mmio_req_bits_size),
    .io_mmio_req_bits_cmd(Cache_1_io_mmio_req_bits_cmd),
    .io_mmio_req_bits_wmask(Cache_1_io_mmio_req_bits_wmask),
    .io_mmio_req_bits_wdata(Cache_1_io_mmio_req_bits_wdata),
    .io_mmio_resp_valid(Cache_1_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(Cache_1_io_mmio_resp_bits_rdata),
    .io_empty(Cache_1_io_empty),
    .mmio(Cache_1_mmio),
    .DISPLAY_ENABLE(Cache_1_DISPLAY_ENABLE)
  );
  assign io_imem_mem_req_valid = Cache_io_out_mem_req_valid; // @[NutCore.scala 153:13]
  assign io_imem_mem_req_bits_addr = Cache_io_out_mem_req_bits_addr; // @[NutCore.scala 153:13]
  assign io_imem_mem_req_bits_cmd = Cache_io_out_mem_req_bits_cmd; // @[NutCore.scala 153:13]
  assign io_imem_mem_req_bits_wdata = Cache_io_out_mem_req_bits_wdata; // @[NutCore.scala 153:13]
  assign io_dmem_mem_req_valid = Cache_1_io_out_mem_req_valid; // @[NutCore.scala 158:13]
  assign io_dmem_mem_req_bits_addr = Cache_1_io_out_mem_req_bits_addr; // @[NutCore.scala 158:13]
  assign io_dmem_mem_req_bits_cmd = Cache_1_io_out_mem_req_bits_cmd; // @[NutCore.scala 158:13]
  assign io_dmem_mem_req_bits_wdata = Cache_1_io_out_mem_req_bits_wdata; // @[NutCore.scala 158:13]
  assign io_dmem_coh_req_ready = Cache_1_io_out_coh_req_ready; // @[NutCore.scala 158:13]
  assign io_dmem_coh_resp_valid = Cache_1_io_out_coh_resp_valid; // @[NutCore.scala 158:13]
  assign io_dmem_coh_resp_bits_cmd = Cache_1_io_out_coh_resp_bits_cmd; // @[NutCore.scala 158:13]
  assign io_dmem_coh_resp_bits_rdata = Cache_1_io_out_coh_resp_bits_rdata; // @[NutCore.scala 158:13]
  assign io_mmio_req_valid = SimpleBusCrossbarNto1_io_out_req_valid; // @[NutCore.scala 167:13]
  assign io_mmio_req_bits_addr = SimpleBusCrossbarNto1_io_out_req_bits_addr; // @[NutCore.scala 167:13]
  assign io_mmio_req_bits_size = SimpleBusCrossbarNto1_io_out_req_bits_size; // @[NutCore.scala 167:13]
  assign io_mmio_req_bits_cmd = SimpleBusCrossbarNto1_io_out_req_bits_cmd; // @[NutCore.scala 167:13]
  assign io_mmio_req_bits_wmask = SimpleBusCrossbarNto1_io_out_req_bits_wmask; // @[NutCore.scala 167:13]
  assign io_mmio_req_bits_wdata = SimpleBusCrossbarNto1_io_out_req_bits_wdata; // @[NutCore.scala 167:13]
  assign io_frontend_req_ready = SimpleBusCrossbarNto1_1_io_in_3_req_ready; // @[NutCore.scala 165:23]
  assign io_frontend_resp_valid = SimpleBusCrossbarNto1_1_io_in_3_resp_valid; // @[NutCore.scala 165:23]
  assign io_frontend_resp_bits_cmd = SimpleBusCrossbarNto1_1_io_in_3_resp_bits_cmd; // @[NutCore.scala 165:23]
  assign io_frontend_resp_bits_rdata = SimpleBusCrossbarNto1_1_io_in_3_resp_bits_rdata; // @[NutCore.scala 165:23]
  assign _T_4181 = Backend_inorder__T_4181;
  assign _T_4184 = Backend_inorder__T_4184;
  assign _T_4185 = Backend_inorder__T_4185;
  assign falseWire = Backend_inorder_falseWire;
  assign falseWire_0 = Backend_inorder_falseWire_0;
  assign _T_4178 = Backend_inorder__T_4178;
  assign _T_284_0 = Backend_inorder__T_284_0;
  assign _T_284_1 = Backend_inorder__T_284_1;
  assign _T_284_2 = Backend_inorder__T_284_2;
  assign _T_284_3 = Backend_inorder__T_284_3;
  assign _T_284_4 = Backend_inorder__T_284_4;
  assign _T_284_5 = Backend_inorder__T_284_5;
  assign _T_284_6 = Backend_inorder__T_284_6;
  assign _T_284_7 = Backend_inorder__T_284_7;
  assign _T_284_8 = Backend_inorder__T_284_8;
  assign _T_284_9 = Backend_inorder__T_284_9;
  assign _T_284_10 = Backend_inorder__T_284_10;
  assign _T_284_11 = Backend_inorder__T_284_11;
  assign _T_284_12 = Backend_inorder__T_284_12;
  assign _T_284_13 = Backend_inorder__T_284_13;
  assign _T_284_14 = Backend_inorder__T_284_14;
  assign _T_284_15 = Backend_inorder__T_284_15;
  assign _T_284_16 = Backend_inorder__T_284_16;
  assign _T_284_17 = Backend_inorder__T_284_17;
  assign _T_284_18 = Backend_inorder__T_284_18;
  assign _T_284_19 = Backend_inorder__T_284_19;
  assign _T_284_20 = Backend_inorder__T_284_20;
  assign _T_284_21 = Backend_inorder__T_284_21;
  assign _T_284_22 = Backend_inorder__T_284_22;
  assign _T_284_23 = Backend_inorder__T_284_23;
  assign _T_284_24 = Backend_inorder__T_284_24;
  assign _T_284_25 = Backend_inorder__T_284_25;
  assign _T_284_26 = Backend_inorder__T_284_26;
  assign _T_284_27 = Backend_inorder__T_284_27;
  assign _T_284_28 = Backend_inorder__T_284_28;
  assign _T_284_29 = Backend_inorder__T_284_29;
  assign _T_284_30 = Backend_inorder__T_284_30;
  assign _T_284_31 = Backend_inorder__T_284_31;
  assign _T_36_0 = Backend_inorder__T_36;
  assign _T_32_0 = Backend_inorder__T_32;
  assign _T_31_0 = Backend_inorder__T_31;
  assign _T_37_0 = Backend_inorder__T_37;
  assign _T_26_0 = Backend_inorder__T_26;
  assign _T_0 = frontend__T_0;
  assign _T_4183 = Backend_inorder__T_4183;
  assign _T_4182 = Backend_inorder__T_4182;
  assign _T_33_0 = Backend_inorder__T_33;
  assign _T_4179 = Backend_inorder__T_4179;
  assign frontend_clock = clock;
  assign frontend_reset = reset;
  assign frontend_io_out_0_ready = _T_17 | _T_32; // @[PipelineVector.scala 50:15]
  assign frontend_io_imem_req_ready = EmbeddedTLB_io_in_req_ready; // @[EmbeddedTLB.scala 428:17]
  assign frontend_io_imem_resp_valid = EmbeddedTLB_io_in_resp_valid; // @[EmbeddedTLB.scala 428:17]
  assign frontend_io_imem_resp_bits_rdata = EmbeddedTLB_io_in_resp_bits_rdata; // @[EmbeddedTLB.scala 428:17]
  assign frontend_io_imem_resp_bits_user = EmbeddedTLB_io_in_resp_bits_user; // @[EmbeddedTLB.scala 428:17]
  assign frontend_io_ipf = EmbeddedTLB_io_ipf; // @[NutCore.scala 152:21]
  assign frontend_io_redirect_target = Backend_inorder_io_redirect_target; // @[NutCore.scala 161:26]
  assign frontend_io_redirect_valid = Backend_inorder_io_redirect_valid; // @[NutCore.scala 161:26]
  assign frontend_flushICache = Backend_inorder_flushICache;
  assign frontend__T_243_valid = Backend_inorder__T_243_valid;
  assign frontend__T_243_pc = Backend_inorder__T_243_pc;
  assign frontend__T_243_isMissPredict = Backend_inorder__T_243_isMissPredict;
  assign frontend__T_243_actualTarget = Backend_inorder__T_243_actualTarget;
  assign frontend__T_243_actualTaken = Backend_inorder__T_243_actualTaken;
  assign frontend__T_243_fuOpType = Backend_inorder__T_243_fuOpType;
  assign frontend__T_243_btbType = Backend_inorder__T_243_btbType;
  assign frontend__T_243_isRVC = Backend_inorder__T_243_isRVC;
  assign frontend_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign frontend_vmEnable = EmbeddedTLB_1_vmEnable_0;
  assign frontend_intrVec = Backend_inorder_intrVec;
  assign frontend_flushTLB = Backend_inorder_flushTLB;
  assign Backend_inorder_clock = clock;
  assign Backend_inorder_reset = reset;
  assign Backend_inorder_io_in_0_valid = _T_7 != _T_8; // @[PipelineVector.scala 56:16]
  assign Backend_inorder_io_in_0_bits_cf_instr = 2'h3 == _T_8 ? _T_6_3_cf_instr : _GEN_1321; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_pc = 2'h3 == _T_8 ? _T_6_3_cf_pc : _GEN_1322; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_pnpc = 2'h3 == _T_8 ? _T_6_3_cf_pnpc : _GEN_1323; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_exceptionVec_1 = 2'h3 == _T_8 ? _T_6_3_cf_exceptionVec_1 : _GEN_1328; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_exceptionVec_2 = 2'h3 == _T_8 ? _T_6_3_cf_exceptionVec_2 : _GEN_1329; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_exceptionVec_12 = 2'h3 == _T_8 ? _T_6_3_cf_exceptionVec_12 : _GEN_1339; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_0 = 2'h3 == _T_8 ? _T_6_3_cf_intrVec_0 : _GEN_1343; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_1 = 2'h3 == _T_8 ? _T_6_3_cf_intrVec_1 : _GEN_1344; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_2 = 2'h3 == _T_8 ? _T_6_3_cf_intrVec_2 : _GEN_1345; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_3 = 2'h3 == _T_8 ? _T_6_3_cf_intrVec_3 : _GEN_1346; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_4 = 2'h3 == _T_8 ? _T_6_3_cf_intrVec_4 : _GEN_1347; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_5 = 2'h3 == _T_8 ? _T_6_3_cf_intrVec_5 : _GEN_1348; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_6 = 2'h3 == _T_8 ? _T_6_3_cf_intrVec_6 : _GEN_1349; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_7 = 2'h3 == _T_8 ? _T_6_3_cf_intrVec_7 : _GEN_1350; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_8 = 2'h3 == _T_8 ? _T_6_3_cf_intrVec_8 : _GEN_1351; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_9 = 2'h3 == _T_8 ? _T_6_3_cf_intrVec_9 : _GEN_1352; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_10 = 2'h3 == _T_8 ? _T_6_3_cf_intrVec_10 : _GEN_1353; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_11 = 2'h3 == _T_8 ? _T_6_3_cf_intrVec_11 : _GEN_1354; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_brIdx = 2'h3 == _T_8 ? _T_6_3_cf_brIdx : _GEN_1355; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_crossPageIPFFix = 2'h3 == _T_8 ? _T_6_3_cf_crossPageIPFFix : _GEN_1357; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_ctrl_src1Type = 2'h3 == _T_8 ? _T_6_3_ctrl_src1Type : _GEN_1358; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_ctrl_src2Type = 2'h3 == _T_8 ? _T_6_3_ctrl_src2Type : _GEN_1359; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_ctrl_fuType = 2'h3 == _T_8 ? _T_6_3_ctrl_fuType : _GEN_1360; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_ctrl_fuOpType = 2'h3 == _T_8 ? _T_6_3_ctrl_fuOpType : _GEN_1361; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_ctrl_rfSrc1 = 2'h3 == _T_8 ? _T_6_3_ctrl_rfSrc1 : _GEN_1362; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_ctrl_rfSrc2 = 2'h3 == _T_8 ? _T_6_3_ctrl_rfSrc2 : _GEN_1363; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_ctrl_rfWen = 2'h3 == _T_8 ? _T_6_3_ctrl_rfWen : _GEN_1364; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_ctrl_rfDest = 2'h3 == _T_8 ? _T_6_3_ctrl_rfDest : _GEN_1365; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_ctrl_isNutCoreTrap = 2'h3 == _T_8 ? _T_6_3_ctrl_isNutCoreTrap : _GEN_1368; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_data_imm = 2'h3 == _T_8 ? _T_6_3_data_imm : _GEN_1375; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_flush = frontend_io_flushVec[3:2]; // @[NutCore.scala 162:22]
  assign Backend_inorder_io_dmem_req_ready = EmbeddedTLB_1_io_in_req_ready; // @[EmbeddedTLB.scala 428:17]
  assign Backend_inorder_io_dmem_resp_valid = EmbeddedTLB_1_io_in_resp_valid; // @[EmbeddedTLB.scala 428:17]
  assign Backend_inorder_io_dmem_resp_bits_rdata = EmbeddedTLB_1_io_in_resp_bits_rdata; // @[EmbeddedTLB.scala 428:17]
  assign Backend_inorder_io_memMMU_dmem_loadPF = EmbeddedTLB_1_io_csrMMU_loadPF; // @[EmbeddedTLB.scala 431:21]
  assign Backend_inorder_io_memMMU_dmem_storePF = EmbeddedTLB_1_io_csrMMU_storePF; // @[EmbeddedTLB.scala 431:21]
  assign Backend_inorder_io_memMMU_dmem_addr = EmbeddedTLB_1_io_csrMMU_addr; // @[EmbeddedTLB.scala 431:21]
  assign Backend_inorder__T_38 = EmbeddedTLB_1__T_38_0;
  assign Backend_inorder_mmio = Cache_1_mmio;
  assign Backend_inorder_io_extra_mtip = io_extra_mtip;
  assign Backend_inorder__T_13 = DISPLAY_ENABLE;
  assign Backend_inorder_io_extra_meip_0 = io_extra_meip_0;
  assign Backend_inorder_vmEnable = EmbeddedTLB_1_vmEnable_0;
  assign Backend_inorder__T_37_0 = EmbeddedTLB_1__T_37_1;
  assign Backend_inorder_io_extra_msip = io_extra_msip;
  assign Backend_inorder__T_65 = frontend__T_65;
  assign Backend_inorder__T_66 = frontend__T_66;
  assign SimpleBusCrossbarNto1_clock = clock;
  assign SimpleBusCrossbarNto1_reset = reset;
  assign SimpleBusCrossbarNto1_io_in_0_req_valid = Cache_io_mmio_req_valid; // @[Cache.scala 685:13]
  assign SimpleBusCrossbarNto1_io_in_0_req_bits_addr = Cache_io_mmio_req_bits_addr; // @[Cache.scala 685:13]
  assign SimpleBusCrossbarNto1_io_in_0_req_bits_cmd = 4'h0; // @[Cache.scala 685:13]
  assign SimpleBusCrossbarNto1_io_in_0_req_bits_wmask = 8'h0; // @[Cache.scala 685:13]
  assign SimpleBusCrossbarNto1_io_in_0_req_bits_wdata = 64'h0; // @[Cache.scala 685:13]
  assign SimpleBusCrossbarNto1_io_in_1_req_valid = Cache_1_io_mmio_req_valid; // @[Cache.scala 685:13]
  assign SimpleBusCrossbarNto1_io_in_1_req_bits_addr = Cache_1_io_mmio_req_bits_addr; // @[Cache.scala 685:13]
  assign SimpleBusCrossbarNto1_io_in_1_req_bits_size = Cache_1_io_mmio_req_bits_size; // @[Cache.scala 685:13]
  assign SimpleBusCrossbarNto1_io_in_1_req_bits_cmd = Cache_1_io_mmio_req_bits_cmd; // @[Cache.scala 685:13]
  assign SimpleBusCrossbarNto1_io_in_1_req_bits_wmask = Cache_1_io_mmio_req_bits_wmask; // @[Cache.scala 685:13]
  assign SimpleBusCrossbarNto1_io_in_1_req_bits_wdata = Cache_1_io_mmio_req_bits_wdata; // @[Cache.scala 685:13]
  assign SimpleBusCrossbarNto1_io_out_req_ready = io_mmio_req_ready; // @[NutCore.scala 167:13]
  assign SimpleBusCrossbarNto1_io_out_resp_valid = io_mmio_resp_valid; // @[NutCore.scala 167:13]
  assign SimpleBusCrossbarNto1_io_out_resp_bits_cmd = 4'h6; // @[NutCore.scala 167:13]
  assign SimpleBusCrossbarNto1_io_out_resp_bits_rdata = io_mmio_resp_bits_rdata; // @[NutCore.scala 167:13]
  assign SimpleBusCrossbarNto1_1_clock = clock;
  assign SimpleBusCrossbarNto1_1_reset = reset;
  assign SimpleBusCrossbarNto1_1_io_in_0_req_valid = EmbeddedTLB_1_io_out_req_valid; // @[NutCore.scala 157:23]
  assign SimpleBusCrossbarNto1_1_io_in_0_req_bits_addr = EmbeddedTLB_1_io_out_req_bits_addr; // @[NutCore.scala 157:23]
  assign SimpleBusCrossbarNto1_1_io_in_0_req_bits_size = EmbeddedTLB_1_io_out_req_bits_size; // @[NutCore.scala 157:23]
  assign SimpleBusCrossbarNto1_1_io_in_0_req_bits_cmd = EmbeddedTLB_1_io_out_req_bits_cmd; // @[NutCore.scala 157:23]
  assign SimpleBusCrossbarNto1_1_io_in_0_req_bits_wmask = EmbeddedTLB_1_io_out_req_bits_wmask; // @[NutCore.scala 157:23]
  assign SimpleBusCrossbarNto1_1_io_in_0_req_bits_wdata = EmbeddedTLB_1_io_out_req_bits_wdata; // @[NutCore.scala 157:23]
  assign SimpleBusCrossbarNto1_1_io_in_1_req_valid = EmbeddedTLB_io_mem_req_valid; // @[EmbeddedTLB.scala 429:18]
  assign SimpleBusCrossbarNto1_1_io_in_1_req_bits_addr = EmbeddedTLB_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 429:18]
  assign SimpleBusCrossbarNto1_1_io_in_1_req_bits_cmd = EmbeddedTLB_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 429:18]
  assign SimpleBusCrossbarNto1_1_io_in_1_req_bits_wdata = EmbeddedTLB_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 429:18]
  assign SimpleBusCrossbarNto1_1_io_in_2_req_valid = EmbeddedTLB_1_io_mem_req_valid; // @[EmbeddedTLB.scala 429:18]
  assign SimpleBusCrossbarNto1_1_io_in_2_req_bits_addr = EmbeddedTLB_1_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 429:18]
  assign SimpleBusCrossbarNto1_1_io_in_2_req_bits_cmd = EmbeddedTLB_1_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 429:18]
  assign SimpleBusCrossbarNto1_1_io_in_2_req_bits_wdata = EmbeddedTLB_1_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 429:18]
  assign SimpleBusCrossbarNto1_1_io_in_3_req_valid = io_frontend_req_valid; // @[NutCore.scala 165:23]
  assign SimpleBusCrossbarNto1_1_io_in_3_req_bits_addr = io_frontend_req_bits_addr; // @[NutCore.scala 165:23]
  assign SimpleBusCrossbarNto1_1_io_in_3_req_bits_size = io_frontend_req_bits_size; // @[NutCore.scala 165:23]
  assign SimpleBusCrossbarNto1_1_io_in_3_req_bits_cmd = io_frontend_req_bits_cmd; // @[NutCore.scala 165:23]
  assign SimpleBusCrossbarNto1_1_io_in_3_req_bits_wmask = io_frontend_req_bits_wmask; // @[NutCore.scala 165:23]
  assign SimpleBusCrossbarNto1_1_io_in_3_req_bits_wdata = io_frontend_req_bits_wdata; // @[NutCore.scala 165:23]
  assign SimpleBusCrossbarNto1_1_io_in_3_resp_ready = io_frontend_resp_ready; // @[NutCore.scala 165:23]
  assign SimpleBusCrossbarNto1_1_io_out_req_ready = Cache_1_io_in_req_ready; // @[Cache.scala 684:17]
  assign SimpleBusCrossbarNto1_1_io_out_resp_valid = Cache_1_io_in_resp_valid; // @[Cache.scala 684:17]
  assign SimpleBusCrossbarNto1_1_io_out_resp_bits_cmd = Cache_1_io_in_resp_bits_cmd; // @[Cache.scala 684:17]
  assign SimpleBusCrossbarNto1_1_io_out_resp_bits_rdata = Cache_1_io_in_resp_bits_rdata; // @[Cache.scala 684:17]
  assign EmbeddedTLB_clock = clock;
  assign EmbeddedTLB_reset = reset;
  assign EmbeddedTLB_io_in_req_valid = frontend_io_imem_req_valid; // @[EmbeddedTLB.scala 428:17]
  assign EmbeddedTLB_io_in_req_bits_addr = frontend_io_imem_req_bits_addr; // @[EmbeddedTLB.scala 428:17]
  assign EmbeddedTLB_io_in_req_bits_user = frontend_io_imem_req_bits_user; // @[EmbeddedTLB.scala 428:17]
  assign EmbeddedTLB_io_in_resp_ready = frontend_io_imem_resp_ready; // @[EmbeddedTLB.scala 428:17]
  assign EmbeddedTLB_io_out_req_ready = Cache_io_in_req_ready; // @[Cache.scala 684:17]
  assign EmbeddedTLB_io_out_resp_valid = Cache_io_in_resp_valid; // @[Cache.scala 684:17]
  assign EmbeddedTLB_io_out_resp_bits_rdata = Cache_io_in_resp_bits_rdata; // @[Cache.scala 684:17]
  assign EmbeddedTLB_io_out_resp_bits_user = Cache_io_in_resp_bits_user; // @[Cache.scala 684:17]
  assign EmbeddedTLB_io_mem_req_ready = SimpleBusCrossbarNto1_1_io_in_1_req_ready; // @[EmbeddedTLB.scala 429:18]
  assign EmbeddedTLB_io_mem_resp_valid = SimpleBusCrossbarNto1_1_io_in_1_resp_valid; // @[EmbeddedTLB.scala 429:18]
  assign EmbeddedTLB_io_mem_resp_bits_cmd = SimpleBusCrossbarNto1_1_io_in_1_resp_bits_cmd; // @[EmbeddedTLB.scala 429:18]
  assign EmbeddedTLB_io_mem_resp_bits_rdata = SimpleBusCrossbarNto1_1_io_in_1_resp_bits_rdata; // @[EmbeddedTLB.scala 429:18]
  assign EmbeddedTLB_io_flush = frontend_io_flushVec[0]; // @[EmbeddedTLB.scala 430:20]
  assign EmbeddedTLB_io_csrMMU_priviledgeMode = Backend_inorder_io_memMMU_imem_priviledgeMode; // @[EmbeddedTLB.scala 431:21]
  assign EmbeddedTLB_io_cacheEmpty = Cache_io_empty; // @[Cache.scala 686:11]
  assign EmbeddedTLB_CSRSATP = Backend_inorder_satp;
  assign EmbeddedTLB_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign EmbeddedTLB_MOUFlushTLB = Backend_inorder_flushTLB;
  assign Cache_clock = clock;
  assign Cache_reset = reset;
  assign Cache_io_in_req_valid = EmbeddedTLB_io_out_req_valid; // @[Cache.scala 684:17]
  assign Cache_io_in_req_bits_addr = EmbeddedTLB_io_out_req_bits_addr; // @[Cache.scala 684:17]
  assign Cache_io_in_req_bits_user = EmbeddedTLB_io_out_req_bits_user; // @[Cache.scala 684:17]
  assign Cache_io_in_resp_ready = EmbeddedTLB_io_out_resp_ready; // @[Cache.scala 684:17]
  assign Cache_io_flush = frontend_io_flushVec[0] ? 2'h3 : 2'h0; // @[Cache.scala 683:20]
  assign Cache_io_out_mem_req_ready = io_imem_mem_req_ready; // @[NutCore.scala 153:13]
  assign Cache_io_out_mem_resp_valid = io_imem_mem_resp_valid; // @[NutCore.scala 153:13]
  assign Cache_io_out_mem_resp_bits_cmd = io_imem_mem_resp_bits_cmd; // @[NutCore.scala 153:13]
  assign Cache_io_out_mem_resp_bits_rdata = io_imem_mem_resp_bits_rdata; // @[NutCore.scala 153:13]
  assign Cache_io_mmio_req_ready = SimpleBusCrossbarNto1_io_in_0_req_ready; // @[Cache.scala 685:13]
  assign Cache_io_mmio_resp_valid = SimpleBusCrossbarNto1_io_in_0_resp_valid; // @[Cache.scala 685:13]
  assign Cache_io_mmio_resp_bits_rdata = SimpleBusCrossbarNto1_io_in_0_resp_bits_rdata; // @[Cache.scala 685:13]
  assign Cache_MOUFlushICache = Backend_inorder_flushICache;
  assign Cache_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign EmbeddedTLB_1_clock = clock;
  assign EmbeddedTLB_1_reset = reset;
  assign EmbeddedTLB_1_io_in_req_valid = Backend_inorder_io_dmem_req_valid; // @[EmbeddedTLB.scala 428:17]
  assign EmbeddedTLB_1_io_in_req_bits_addr = Backend_inorder_io_dmem_req_bits_addr; // @[EmbeddedTLB.scala 428:17]
  assign EmbeddedTLB_1_io_in_req_bits_size = Backend_inorder_io_dmem_req_bits_size; // @[EmbeddedTLB.scala 428:17]
  assign EmbeddedTLB_1_io_in_req_bits_cmd = Backend_inorder_io_dmem_req_bits_cmd; // @[EmbeddedTLB.scala 428:17]
  assign EmbeddedTLB_1_io_in_req_bits_wmask = Backend_inorder_io_dmem_req_bits_wmask; // @[EmbeddedTLB.scala 428:17]
  assign EmbeddedTLB_1_io_in_req_bits_wdata = Backend_inorder_io_dmem_req_bits_wdata; // @[EmbeddedTLB.scala 428:17]
  assign EmbeddedTLB_1_io_out_req_ready = SimpleBusCrossbarNto1_1_io_in_0_req_ready; // @[NutCore.scala 157:23]
  assign EmbeddedTLB_1_io_out_resp_valid = SimpleBusCrossbarNto1_1_io_in_0_resp_valid; // @[NutCore.scala 157:23]
  assign EmbeddedTLB_1_io_out_resp_bits_cmd = SimpleBusCrossbarNto1_1_io_in_0_resp_bits_cmd; // @[NutCore.scala 157:23]
  assign EmbeddedTLB_1_io_out_resp_bits_rdata = SimpleBusCrossbarNto1_1_io_in_0_resp_bits_rdata; // @[NutCore.scala 157:23]
  assign EmbeddedTLB_1_io_mem_req_ready = SimpleBusCrossbarNto1_1_io_in_2_req_ready; // @[EmbeddedTLB.scala 429:18]
  assign EmbeddedTLB_1_io_mem_resp_valid = SimpleBusCrossbarNto1_1_io_in_2_resp_valid; // @[EmbeddedTLB.scala 429:18]
  assign EmbeddedTLB_1_io_mem_resp_bits_cmd = SimpleBusCrossbarNto1_1_io_in_2_resp_bits_cmd; // @[EmbeddedTLB.scala 429:18]
  assign EmbeddedTLB_1_io_mem_resp_bits_rdata = SimpleBusCrossbarNto1_1_io_in_2_resp_bits_rdata; // @[EmbeddedTLB.scala 429:18]
  assign EmbeddedTLB_1_io_csrMMU_priviledgeMode = Backend_inorder_io_memMMU_dmem_priviledgeMode; // @[EmbeddedTLB.scala 431:21]
  assign EmbeddedTLB_1_io_csrMMU_status_sum = Backend_inorder_io_memMMU_dmem_status_sum; // @[EmbeddedTLB.scala 431:21]
  assign EmbeddedTLB_1_io_csrMMU_status_mxr = Backend_inorder_io_memMMU_dmem_status_mxr; // @[EmbeddedTLB.scala 431:21]
  assign EmbeddedTLB_1_io_cacheEmpty = Cache_1_io_empty; // @[Cache.scala 686:11]
  assign EmbeddedTLB_1_CSRSATP = Backend_inorder_satp;
  assign EmbeddedTLB_1_amoReq = Backend_inorder_amoReq;
  assign EmbeddedTLB_1_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign EmbeddedTLB_1_MOUFlushTLB = Backend_inorder_flushTLB;
  assign Cache_1_clock = clock;
  assign Cache_1_reset = reset;
  assign Cache_1_io_in_req_valid = SimpleBusCrossbarNto1_1_io_out_req_valid; // @[Cache.scala 684:17]
  assign Cache_1_io_in_req_bits_addr = SimpleBusCrossbarNto1_1_io_out_req_bits_addr; // @[Cache.scala 684:17]
  assign Cache_1_io_in_req_bits_size = SimpleBusCrossbarNto1_1_io_out_req_bits_size; // @[Cache.scala 684:17]
  assign Cache_1_io_in_req_bits_cmd = SimpleBusCrossbarNto1_1_io_out_req_bits_cmd; // @[Cache.scala 684:17]
  assign Cache_1_io_in_req_bits_wmask = SimpleBusCrossbarNto1_1_io_out_req_bits_wmask; // @[Cache.scala 684:17]
  assign Cache_1_io_in_req_bits_wdata = SimpleBusCrossbarNto1_1_io_out_req_bits_wdata; // @[Cache.scala 684:17]
  assign Cache_1_io_in_resp_ready = SimpleBusCrossbarNto1_1_io_out_resp_ready; // @[Cache.scala 684:17]
  assign Cache_1_io_out_mem_req_ready = io_dmem_mem_req_ready; // @[NutCore.scala 158:13]
  assign Cache_1_io_out_mem_resp_valid = io_dmem_mem_resp_valid; // @[NutCore.scala 158:13]
  assign Cache_1_io_out_mem_resp_bits_cmd = io_dmem_mem_resp_bits_cmd; // @[NutCore.scala 158:13]
  assign Cache_1_io_out_mem_resp_bits_rdata = io_dmem_mem_resp_bits_rdata; // @[NutCore.scala 158:13]
  assign Cache_1_io_out_coh_req_valid = io_dmem_coh_req_valid; // @[NutCore.scala 158:13]
  assign Cache_1_io_out_coh_req_bits_addr = io_dmem_coh_req_bits_addr; // @[NutCore.scala 158:13]
  assign Cache_1_io_out_coh_req_bits_wdata = io_dmem_coh_req_bits_wdata; // @[NutCore.scala 158:13]
  assign Cache_1_io_mmio_req_ready = SimpleBusCrossbarNto1_io_in_1_req_ready; // @[Cache.scala 685:13]
  assign Cache_1_io_mmio_resp_valid = SimpleBusCrossbarNto1_io_in_1_resp_valid; // @[Cache.scala 685:13]
  assign Cache_1_io_mmio_resp_bits_rdata = SimpleBusCrossbarNto1_io_in_1_resp_bits_rdata; // @[Cache.scala 685:13]
  assign Cache_1_DISPLAY_ENABLE = DISPLAY_ENABLE;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  _T_6_0_cf_instr = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  _T_6_0_cf_pc = _RAND_1[38:0];
  _RAND_2 = {2{`RANDOM}};
  _T_6_0_cf_pnpc = _RAND_2[38:0];
  _RAND_3 = {1{`RANDOM}};
  _T_6_0_cf_exceptionVec_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_6_0_cf_exceptionVec_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _T_6_0_cf_exceptionVec_12 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _T_6_0_cf_intrVec_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_6_0_cf_intrVec_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _T_6_0_cf_intrVec_2 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _T_6_0_cf_intrVec_3 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _T_6_0_cf_intrVec_4 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _T_6_0_cf_intrVec_5 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _T_6_0_cf_intrVec_6 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _T_6_0_cf_intrVec_7 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  _T_6_0_cf_intrVec_8 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  _T_6_0_cf_intrVec_9 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  _T_6_0_cf_intrVec_10 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  _T_6_0_cf_intrVec_11 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  _T_6_0_cf_brIdx = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  _T_6_0_cf_crossPageIPFFix = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  _T_6_0_ctrl_src1Type = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  _T_6_0_ctrl_src2Type = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  _T_6_0_ctrl_fuType = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  _T_6_0_ctrl_fuOpType = _RAND_23[6:0];
  _RAND_24 = {1{`RANDOM}};
  _T_6_0_ctrl_rfSrc1 = _RAND_24[4:0];
  _RAND_25 = {1{`RANDOM}};
  _T_6_0_ctrl_rfSrc2 = _RAND_25[4:0];
  _RAND_26 = {1{`RANDOM}};
  _T_6_0_ctrl_rfWen = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  _T_6_0_ctrl_rfDest = _RAND_27[4:0];
  _RAND_28 = {1{`RANDOM}};
  _T_6_0_ctrl_isNutCoreTrap = _RAND_28[0:0];
  _RAND_29 = {2{`RANDOM}};
  _T_6_0_data_imm = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  _T_6_1_cf_instr = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  _T_6_1_cf_pc = _RAND_31[38:0];
  _RAND_32 = {2{`RANDOM}};
  _T_6_1_cf_pnpc = _RAND_32[38:0];
  _RAND_33 = {1{`RANDOM}};
  _T_6_1_cf_exceptionVec_1 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  _T_6_1_cf_exceptionVec_2 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  _T_6_1_cf_exceptionVec_12 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  _T_6_1_cf_intrVec_0 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  _T_6_1_cf_intrVec_1 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  _T_6_1_cf_intrVec_2 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  _T_6_1_cf_intrVec_3 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  _T_6_1_cf_intrVec_4 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  _T_6_1_cf_intrVec_5 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  _T_6_1_cf_intrVec_6 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  _T_6_1_cf_intrVec_7 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  _T_6_1_cf_intrVec_8 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  _T_6_1_cf_intrVec_9 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  _T_6_1_cf_intrVec_10 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  _T_6_1_cf_intrVec_11 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  _T_6_1_cf_brIdx = _RAND_48[3:0];
  _RAND_49 = {1{`RANDOM}};
  _T_6_1_cf_crossPageIPFFix = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  _T_6_1_ctrl_src1Type = _RAND_50[1:0];
  _RAND_51 = {1{`RANDOM}};
  _T_6_1_ctrl_src2Type = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  _T_6_1_ctrl_fuType = _RAND_52[2:0];
  _RAND_53 = {1{`RANDOM}};
  _T_6_1_ctrl_fuOpType = _RAND_53[6:0];
  _RAND_54 = {1{`RANDOM}};
  _T_6_1_ctrl_rfSrc1 = _RAND_54[4:0];
  _RAND_55 = {1{`RANDOM}};
  _T_6_1_ctrl_rfSrc2 = _RAND_55[4:0];
  _RAND_56 = {1{`RANDOM}};
  _T_6_1_ctrl_rfWen = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  _T_6_1_ctrl_rfDest = _RAND_57[4:0];
  _RAND_58 = {1{`RANDOM}};
  _T_6_1_ctrl_isNutCoreTrap = _RAND_58[0:0];
  _RAND_59 = {2{`RANDOM}};
  _T_6_1_data_imm = _RAND_59[63:0];
  _RAND_60 = {2{`RANDOM}};
  _T_6_2_cf_instr = _RAND_60[63:0];
  _RAND_61 = {2{`RANDOM}};
  _T_6_2_cf_pc = _RAND_61[38:0];
  _RAND_62 = {2{`RANDOM}};
  _T_6_2_cf_pnpc = _RAND_62[38:0];
  _RAND_63 = {1{`RANDOM}};
  _T_6_2_cf_exceptionVec_1 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  _T_6_2_cf_exceptionVec_2 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  _T_6_2_cf_exceptionVec_12 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  _T_6_2_cf_intrVec_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  _T_6_2_cf_intrVec_1 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  _T_6_2_cf_intrVec_2 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  _T_6_2_cf_intrVec_3 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  _T_6_2_cf_intrVec_4 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  _T_6_2_cf_intrVec_5 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  _T_6_2_cf_intrVec_6 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  _T_6_2_cf_intrVec_7 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  _T_6_2_cf_intrVec_8 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  _T_6_2_cf_intrVec_9 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  _T_6_2_cf_intrVec_10 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  _T_6_2_cf_intrVec_11 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  _T_6_2_cf_brIdx = _RAND_78[3:0];
  _RAND_79 = {1{`RANDOM}};
  _T_6_2_cf_crossPageIPFFix = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  _T_6_2_ctrl_src1Type = _RAND_80[1:0];
  _RAND_81 = {1{`RANDOM}};
  _T_6_2_ctrl_src2Type = _RAND_81[1:0];
  _RAND_82 = {1{`RANDOM}};
  _T_6_2_ctrl_fuType = _RAND_82[2:0];
  _RAND_83 = {1{`RANDOM}};
  _T_6_2_ctrl_fuOpType = _RAND_83[6:0];
  _RAND_84 = {1{`RANDOM}};
  _T_6_2_ctrl_rfSrc1 = _RAND_84[4:0];
  _RAND_85 = {1{`RANDOM}};
  _T_6_2_ctrl_rfSrc2 = _RAND_85[4:0];
  _RAND_86 = {1{`RANDOM}};
  _T_6_2_ctrl_rfWen = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  _T_6_2_ctrl_rfDest = _RAND_87[4:0];
  _RAND_88 = {1{`RANDOM}};
  _T_6_2_ctrl_isNutCoreTrap = _RAND_88[0:0];
  _RAND_89 = {2{`RANDOM}};
  _T_6_2_data_imm = _RAND_89[63:0];
  _RAND_90 = {2{`RANDOM}};
  _T_6_3_cf_instr = _RAND_90[63:0];
  _RAND_91 = {2{`RANDOM}};
  _T_6_3_cf_pc = _RAND_91[38:0];
  _RAND_92 = {2{`RANDOM}};
  _T_6_3_cf_pnpc = _RAND_92[38:0];
  _RAND_93 = {1{`RANDOM}};
  _T_6_3_cf_exceptionVec_1 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  _T_6_3_cf_exceptionVec_2 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  _T_6_3_cf_exceptionVec_12 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  _T_6_3_cf_intrVec_0 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  _T_6_3_cf_intrVec_1 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  _T_6_3_cf_intrVec_2 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  _T_6_3_cf_intrVec_3 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  _T_6_3_cf_intrVec_4 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  _T_6_3_cf_intrVec_5 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  _T_6_3_cf_intrVec_6 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  _T_6_3_cf_intrVec_7 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  _T_6_3_cf_intrVec_8 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  _T_6_3_cf_intrVec_9 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  _T_6_3_cf_intrVec_10 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  _T_6_3_cf_intrVec_11 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  _T_6_3_cf_brIdx = _RAND_108[3:0];
  _RAND_109 = {1{`RANDOM}};
  _T_6_3_cf_crossPageIPFFix = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  _T_6_3_ctrl_src1Type = _RAND_110[1:0];
  _RAND_111 = {1{`RANDOM}};
  _T_6_3_ctrl_src2Type = _RAND_111[1:0];
  _RAND_112 = {1{`RANDOM}};
  _T_6_3_ctrl_fuType = _RAND_112[2:0];
  _RAND_113 = {1{`RANDOM}};
  _T_6_3_ctrl_fuOpType = _RAND_113[6:0];
  _RAND_114 = {1{`RANDOM}};
  _T_6_3_ctrl_rfSrc1 = _RAND_114[4:0];
  _RAND_115 = {1{`RANDOM}};
  _T_6_3_ctrl_rfSrc2 = _RAND_115[4:0];
  _RAND_116 = {1{`RANDOM}};
  _T_6_3_ctrl_rfWen = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  _T_6_3_ctrl_rfDest = _RAND_117[4:0];
  _RAND_118 = {1{`RANDOM}};
  _T_6_3_ctrl_isNutCoreTrap = _RAND_118[0:0];
  _RAND_119 = {2{`RANDOM}};
  _T_6_3_data_imm = _RAND_119[63:0];
  _RAND_120 = {1{`RANDOM}};
  _T_7 = _RAND_120[1:0];
  _RAND_121 = {1{`RANDOM}};
  _T_8 = _RAND_121[1:0];
  _RAND_122 = {2{`RANDOM}};
  _T_62 = _RAND_122[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_6_0_cf_instr <= 64'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_instr <= 64'h0;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_cf_instr <= frontend_io_out_0_bits_cf_instr;
            end else begin
              _T_6_0_cf_instr <= 64'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_cf_instr <= frontend_io_out_0_bits_cf_instr;
          end else begin
            _T_6_0_cf_instr <= 64'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_pc <= 39'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_pc <= 39'h0;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_cf_pc <= frontend_io_out_0_bits_cf_pc;
            end else begin
              _T_6_0_cf_pc <= 39'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_cf_pc <= frontend_io_out_0_bits_cf_pc;
          end else begin
            _T_6_0_cf_pc <= 39'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_pnpc <= 39'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_pnpc <= 39'h0;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_cf_pnpc <= frontend_io_out_0_bits_cf_pnpc;
            end else begin
              _T_6_0_cf_pnpc <= 39'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_cf_pnpc <= frontend_io_out_0_bits_cf_pnpc;
          end else begin
            _T_6_0_cf_pnpc <= 39'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_exceptionVec_1 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_exceptionVec_1 <= 1'h0;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            _T_6_0_cf_exceptionVec_1 <= _T_27_cf_exceptionVec_1;
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          _T_6_0_cf_exceptionVec_1 <= _T_27_cf_exceptionVec_1;
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_exceptionVec_2 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_exceptionVec_2 <= 1'h0;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            _T_6_0_cf_exceptionVec_2 <= _T_27_cf_exceptionVec_2;
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          _T_6_0_cf_exceptionVec_2 <= _T_27_cf_exceptionVec_2;
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_exceptionVec_12 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_exceptionVec_12 <= 1'h0;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            _T_6_0_cf_exceptionVec_12 <= _T_27_cf_exceptionVec_12;
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          _T_6_0_cf_exceptionVec_12 <= _T_27_cf_exceptionVec_12;
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_intrVec_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_intrVec_0 <= _T_6_T_29_cf_intrVec_0;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_cf_intrVec_0 <= frontend_io_out_0_bits_cf_intrVec_0;
            end else begin
              _T_6_0_cf_intrVec_0 <= frontend_io_out_1_bits_cf_intrVec_0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_cf_intrVec_0 <= frontend_io_out_0_bits_cf_intrVec_0;
          end else begin
            _T_6_0_cf_intrVec_0 <= frontend_io_out_1_bits_cf_intrVec_0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_intrVec_1 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_intrVec_1 <= _T_6_T_29_cf_intrVec_1;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_cf_intrVec_1 <= frontend_io_out_0_bits_cf_intrVec_1;
            end else begin
              _T_6_0_cf_intrVec_1 <= frontend_io_out_1_bits_cf_intrVec_1;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_cf_intrVec_1 <= frontend_io_out_0_bits_cf_intrVec_1;
          end else begin
            _T_6_0_cf_intrVec_1 <= frontend_io_out_1_bits_cf_intrVec_1;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_intrVec_2 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_intrVec_2 <= _T_6_T_29_cf_intrVec_2;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_cf_intrVec_2 <= frontend_io_out_0_bits_cf_intrVec_2;
            end else begin
              _T_6_0_cf_intrVec_2 <= frontend_io_out_1_bits_cf_intrVec_2;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_cf_intrVec_2 <= frontend_io_out_0_bits_cf_intrVec_2;
          end else begin
            _T_6_0_cf_intrVec_2 <= frontend_io_out_1_bits_cf_intrVec_2;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_intrVec_3 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_intrVec_3 <= _T_6_T_29_cf_intrVec_3;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_cf_intrVec_3 <= frontend_io_out_0_bits_cf_intrVec_3;
            end else begin
              _T_6_0_cf_intrVec_3 <= frontend_io_out_1_bits_cf_intrVec_3;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_cf_intrVec_3 <= frontend_io_out_0_bits_cf_intrVec_3;
          end else begin
            _T_6_0_cf_intrVec_3 <= frontend_io_out_1_bits_cf_intrVec_3;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_intrVec_4 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_intrVec_4 <= _T_6_T_29_cf_intrVec_4;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_cf_intrVec_4 <= frontend_io_out_0_bits_cf_intrVec_4;
            end else begin
              _T_6_0_cf_intrVec_4 <= frontend_io_out_1_bits_cf_intrVec_4;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_cf_intrVec_4 <= frontend_io_out_0_bits_cf_intrVec_4;
          end else begin
            _T_6_0_cf_intrVec_4 <= frontend_io_out_1_bits_cf_intrVec_4;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_intrVec_5 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_intrVec_5 <= _T_6_T_29_cf_intrVec_5;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_cf_intrVec_5 <= frontend_io_out_0_bits_cf_intrVec_5;
            end else begin
              _T_6_0_cf_intrVec_5 <= frontend_io_out_1_bits_cf_intrVec_5;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_cf_intrVec_5 <= frontend_io_out_0_bits_cf_intrVec_5;
          end else begin
            _T_6_0_cf_intrVec_5 <= frontend_io_out_1_bits_cf_intrVec_5;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_intrVec_6 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_intrVec_6 <= _T_6_T_29_cf_intrVec_6;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_cf_intrVec_6 <= frontend_io_out_0_bits_cf_intrVec_6;
            end else begin
              _T_6_0_cf_intrVec_6 <= frontend_io_out_1_bits_cf_intrVec_6;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_cf_intrVec_6 <= frontend_io_out_0_bits_cf_intrVec_6;
          end else begin
            _T_6_0_cf_intrVec_6 <= frontend_io_out_1_bits_cf_intrVec_6;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_intrVec_7 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_intrVec_7 <= _T_6_T_29_cf_intrVec_7;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_cf_intrVec_7 <= frontend_io_out_0_bits_cf_intrVec_7;
            end else begin
              _T_6_0_cf_intrVec_7 <= frontend_io_out_1_bits_cf_intrVec_7;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_cf_intrVec_7 <= frontend_io_out_0_bits_cf_intrVec_7;
          end else begin
            _T_6_0_cf_intrVec_7 <= frontend_io_out_1_bits_cf_intrVec_7;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_intrVec_8 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_intrVec_8 <= _T_6_T_29_cf_intrVec_8;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_cf_intrVec_8 <= frontend_io_out_0_bits_cf_intrVec_8;
            end else begin
              _T_6_0_cf_intrVec_8 <= frontend_io_out_1_bits_cf_intrVec_8;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_cf_intrVec_8 <= frontend_io_out_0_bits_cf_intrVec_8;
          end else begin
            _T_6_0_cf_intrVec_8 <= frontend_io_out_1_bits_cf_intrVec_8;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_intrVec_9 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_intrVec_9 <= _T_6_T_29_cf_intrVec_9;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_cf_intrVec_9 <= frontend_io_out_0_bits_cf_intrVec_9;
            end else begin
              _T_6_0_cf_intrVec_9 <= frontend_io_out_1_bits_cf_intrVec_9;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_cf_intrVec_9 <= frontend_io_out_0_bits_cf_intrVec_9;
          end else begin
            _T_6_0_cf_intrVec_9 <= frontend_io_out_1_bits_cf_intrVec_9;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_intrVec_10 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_intrVec_10 <= _T_6_T_29_cf_intrVec_10;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_cf_intrVec_10 <= frontend_io_out_0_bits_cf_intrVec_10;
            end else begin
              _T_6_0_cf_intrVec_10 <= frontend_io_out_1_bits_cf_intrVec_10;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_cf_intrVec_10 <= frontend_io_out_0_bits_cf_intrVec_10;
          end else begin
            _T_6_0_cf_intrVec_10 <= frontend_io_out_1_bits_cf_intrVec_10;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_intrVec_11 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_intrVec_11 <= _T_6_T_29_cf_intrVec_11;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_cf_intrVec_11 <= frontend_io_out_0_bits_cf_intrVec_11;
            end else begin
              _T_6_0_cf_intrVec_11 <= frontend_io_out_1_bits_cf_intrVec_11;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_cf_intrVec_11 <= frontend_io_out_0_bits_cf_intrVec_11;
          end else begin
            _T_6_0_cf_intrVec_11 <= frontend_io_out_1_bits_cf_intrVec_11;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_brIdx <= 4'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_brIdx <= 4'h0;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_cf_brIdx <= frontend_io_out_0_bits_cf_brIdx;
            end else begin
              _T_6_0_cf_brIdx <= 4'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_cf_brIdx <= frontend_io_out_0_bits_cf_brIdx;
          end else begin
            _T_6_0_cf_brIdx <= 4'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_crossPageIPFFix <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_crossPageIPFFix <= 1'h0;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            _T_6_0_cf_crossPageIPFFix <= _T_27_cf_crossPageIPFFix;
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          _T_6_0_cf_crossPageIPFFix <= _T_27_cf_crossPageIPFFix;
        end
      end
    end
    if (reset) begin
      _T_6_0_ctrl_src1Type <= 2'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_ctrl_src1Type <= 2'h1;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_ctrl_src1Type <= frontend_io_out_0_bits_ctrl_src1Type;
            end else begin
              _T_6_0_ctrl_src1Type <= 2'h1;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_ctrl_src1Type <= frontend_io_out_0_bits_ctrl_src1Type;
          end else begin
            _T_6_0_ctrl_src1Type <= 2'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_ctrl_src2Type <= 2'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_ctrl_src2Type <= 2'h1;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_ctrl_src2Type <= frontend_io_out_0_bits_ctrl_src2Type;
            end else begin
              _T_6_0_ctrl_src2Type <= 2'h1;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_ctrl_src2Type <= frontend_io_out_0_bits_ctrl_src2Type;
          end else begin
            _T_6_0_ctrl_src2Type <= 2'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_ctrl_fuType <= 3'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_ctrl_fuType <= 3'h3;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_ctrl_fuType <= frontend_io_out_0_bits_ctrl_fuType;
            end else begin
              _T_6_0_ctrl_fuType <= 3'h3;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_ctrl_fuType <= frontend_io_out_0_bits_ctrl_fuType;
          end else begin
            _T_6_0_ctrl_fuType <= 3'h3;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_ctrl_fuOpType <= 7'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_ctrl_fuOpType <= 7'h0;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_ctrl_fuOpType <= frontend_io_out_0_bits_ctrl_fuOpType;
            end else begin
              _T_6_0_ctrl_fuOpType <= 7'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_ctrl_fuOpType <= frontend_io_out_0_bits_ctrl_fuOpType;
          end else begin
            _T_6_0_ctrl_fuOpType <= 7'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_ctrl_rfSrc1 <= 5'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_ctrl_rfSrc1 <= 5'h0;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_ctrl_rfSrc1 <= frontend_io_out_0_bits_ctrl_rfSrc1;
            end else begin
              _T_6_0_ctrl_rfSrc1 <= 5'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_ctrl_rfSrc1 <= frontend_io_out_0_bits_ctrl_rfSrc1;
          end else begin
            _T_6_0_ctrl_rfSrc1 <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_ctrl_rfSrc2 <= 5'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_ctrl_rfSrc2 <= 5'h0;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_ctrl_rfSrc2 <= frontend_io_out_0_bits_ctrl_rfSrc2;
            end else begin
              _T_6_0_ctrl_rfSrc2 <= 5'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_ctrl_rfSrc2 <= frontend_io_out_0_bits_ctrl_rfSrc2;
          end else begin
            _T_6_0_ctrl_rfSrc2 <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_ctrl_rfWen <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_ctrl_rfWen <= 1'h0;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            _T_6_0_ctrl_rfWen <= _T_27_ctrl_rfWen;
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          _T_6_0_ctrl_rfWen <= _T_27_ctrl_rfWen;
        end
      end
    end
    if (reset) begin
      _T_6_0_ctrl_rfDest <= 5'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_ctrl_rfDest <= 5'h0;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_ctrl_rfDest <= frontend_io_out_0_bits_ctrl_rfDest;
            end else begin
              _T_6_0_ctrl_rfDest <= 5'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_ctrl_rfDest <= frontend_io_out_0_bits_ctrl_rfDest;
          end else begin
            _T_6_0_ctrl_rfDest <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_ctrl_isNutCoreTrap <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_ctrl_isNutCoreTrap <= 1'h0;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            _T_6_0_ctrl_isNutCoreTrap <= _T_27_ctrl_isNutCoreTrap;
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          _T_6_0_ctrl_isNutCoreTrap <= _T_27_ctrl_isNutCoreTrap;
        end
      end
    end
    if (reset) begin
      _T_6_0_data_imm <= 64'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_data_imm <= 64'h0;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_data_imm <= frontend_io_out_0_bits_data_imm;
            end else begin
              _T_6_0_data_imm <= 64'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_data_imm <= frontend_io_out_0_bits_data_imm;
          end else begin
            _T_6_0_data_imm <= 64'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_instr <= 64'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_instr <= 64'h0;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_cf_instr <= frontend_io_out_0_bits_cf_instr;
            end else begin
              _T_6_1_cf_instr <= 64'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_cf_instr <= frontend_io_out_0_bits_cf_instr;
          end else begin
            _T_6_1_cf_instr <= 64'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_pc <= 39'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_pc <= 39'h0;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_cf_pc <= frontend_io_out_0_bits_cf_pc;
            end else begin
              _T_6_1_cf_pc <= 39'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_cf_pc <= frontend_io_out_0_bits_cf_pc;
          end else begin
            _T_6_1_cf_pc <= 39'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_pnpc <= 39'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_pnpc <= 39'h0;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_cf_pnpc <= frontend_io_out_0_bits_cf_pnpc;
            end else begin
              _T_6_1_cf_pnpc <= 39'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_cf_pnpc <= frontend_io_out_0_bits_cf_pnpc;
          end else begin
            _T_6_1_cf_pnpc <= 39'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_exceptionVec_1 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_exceptionVec_1 <= 1'h0;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            _T_6_1_cf_exceptionVec_1 <= _T_27_cf_exceptionVec_1;
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          _T_6_1_cf_exceptionVec_1 <= _T_27_cf_exceptionVec_1;
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_exceptionVec_2 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_exceptionVec_2 <= 1'h0;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            _T_6_1_cf_exceptionVec_2 <= _T_27_cf_exceptionVec_2;
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          _T_6_1_cf_exceptionVec_2 <= _T_27_cf_exceptionVec_2;
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_exceptionVec_12 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_exceptionVec_12 <= 1'h0;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            _T_6_1_cf_exceptionVec_12 <= _T_27_cf_exceptionVec_12;
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          _T_6_1_cf_exceptionVec_12 <= _T_27_cf_exceptionVec_12;
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_intrVec_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_intrVec_0 <= _T_6_T_29_cf_intrVec_0;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_cf_intrVec_0 <= frontend_io_out_0_bits_cf_intrVec_0;
            end else begin
              _T_6_1_cf_intrVec_0 <= frontend_io_out_1_bits_cf_intrVec_0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_cf_intrVec_0 <= frontend_io_out_0_bits_cf_intrVec_0;
          end else begin
            _T_6_1_cf_intrVec_0 <= frontend_io_out_1_bits_cf_intrVec_0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_intrVec_1 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_intrVec_1 <= _T_6_T_29_cf_intrVec_1;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_cf_intrVec_1 <= frontend_io_out_0_bits_cf_intrVec_1;
            end else begin
              _T_6_1_cf_intrVec_1 <= frontend_io_out_1_bits_cf_intrVec_1;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_cf_intrVec_1 <= frontend_io_out_0_bits_cf_intrVec_1;
          end else begin
            _T_6_1_cf_intrVec_1 <= frontend_io_out_1_bits_cf_intrVec_1;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_intrVec_2 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_intrVec_2 <= _T_6_T_29_cf_intrVec_2;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_cf_intrVec_2 <= frontend_io_out_0_bits_cf_intrVec_2;
            end else begin
              _T_6_1_cf_intrVec_2 <= frontend_io_out_1_bits_cf_intrVec_2;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_cf_intrVec_2 <= frontend_io_out_0_bits_cf_intrVec_2;
          end else begin
            _T_6_1_cf_intrVec_2 <= frontend_io_out_1_bits_cf_intrVec_2;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_intrVec_3 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_intrVec_3 <= _T_6_T_29_cf_intrVec_3;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_cf_intrVec_3 <= frontend_io_out_0_bits_cf_intrVec_3;
            end else begin
              _T_6_1_cf_intrVec_3 <= frontend_io_out_1_bits_cf_intrVec_3;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_cf_intrVec_3 <= frontend_io_out_0_bits_cf_intrVec_3;
          end else begin
            _T_6_1_cf_intrVec_3 <= frontend_io_out_1_bits_cf_intrVec_3;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_intrVec_4 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_intrVec_4 <= _T_6_T_29_cf_intrVec_4;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_cf_intrVec_4 <= frontend_io_out_0_bits_cf_intrVec_4;
            end else begin
              _T_6_1_cf_intrVec_4 <= frontend_io_out_1_bits_cf_intrVec_4;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_cf_intrVec_4 <= frontend_io_out_0_bits_cf_intrVec_4;
          end else begin
            _T_6_1_cf_intrVec_4 <= frontend_io_out_1_bits_cf_intrVec_4;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_intrVec_5 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_intrVec_5 <= _T_6_T_29_cf_intrVec_5;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_cf_intrVec_5 <= frontend_io_out_0_bits_cf_intrVec_5;
            end else begin
              _T_6_1_cf_intrVec_5 <= frontend_io_out_1_bits_cf_intrVec_5;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_cf_intrVec_5 <= frontend_io_out_0_bits_cf_intrVec_5;
          end else begin
            _T_6_1_cf_intrVec_5 <= frontend_io_out_1_bits_cf_intrVec_5;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_intrVec_6 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_intrVec_6 <= _T_6_T_29_cf_intrVec_6;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_cf_intrVec_6 <= frontend_io_out_0_bits_cf_intrVec_6;
            end else begin
              _T_6_1_cf_intrVec_6 <= frontend_io_out_1_bits_cf_intrVec_6;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_cf_intrVec_6 <= frontend_io_out_0_bits_cf_intrVec_6;
          end else begin
            _T_6_1_cf_intrVec_6 <= frontend_io_out_1_bits_cf_intrVec_6;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_intrVec_7 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_intrVec_7 <= _T_6_T_29_cf_intrVec_7;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_cf_intrVec_7 <= frontend_io_out_0_bits_cf_intrVec_7;
            end else begin
              _T_6_1_cf_intrVec_7 <= frontend_io_out_1_bits_cf_intrVec_7;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_cf_intrVec_7 <= frontend_io_out_0_bits_cf_intrVec_7;
          end else begin
            _T_6_1_cf_intrVec_7 <= frontend_io_out_1_bits_cf_intrVec_7;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_intrVec_8 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_intrVec_8 <= _T_6_T_29_cf_intrVec_8;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_cf_intrVec_8 <= frontend_io_out_0_bits_cf_intrVec_8;
            end else begin
              _T_6_1_cf_intrVec_8 <= frontend_io_out_1_bits_cf_intrVec_8;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_cf_intrVec_8 <= frontend_io_out_0_bits_cf_intrVec_8;
          end else begin
            _T_6_1_cf_intrVec_8 <= frontend_io_out_1_bits_cf_intrVec_8;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_intrVec_9 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_intrVec_9 <= _T_6_T_29_cf_intrVec_9;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_cf_intrVec_9 <= frontend_io_out_0_bits_cf_intrVec_9;
            end else begin
              _T_6_1_cf_intrVec_9 <= frontend_io_out_1_bits_cf_intrVec_9;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_cf_intrVec_9 <= frontend_io_out_0_bits_cf_intrVec_9;
          end else begin
            _T_6_1_cf_intrVec_9 <= frontend_io_out_1_bits_cf_intrVec_9;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_intrVec_10 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_intrVec_10 <= _T_6_T_29_cf_intrVec_10;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_cf_intrVec_10 <= frontend_io_out_0_bits_cf_intrVec_10;
            end else begin
              _T_6_1_cf_intrVec_10 <= frontend_io_out_1_bits_cf_intrVec_10;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_cf_intrVec_10 <= frontend_io_out_0_bits_cf_intrVec_10;
          end else begin
            _T_6_1_cf_intrVec_10 <= frontend_io_out_1_bits_cf_intrVec_10;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_intrVec_11 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_intrVec_11 <= _T_6_T_29_cf_intrVec_11;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_cf_intrVec_11 <= frontend_io_out_0_bits_cf_intrVec_11;
            end else begin
              _T_6_1_cf_intrVec_11 <= frontend_io_out_1_bits_cf_intrVec_11;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_cf_intrVec_11 <= frontend_io_out_0_bits_cf_intrVec_11;
          end else begin
            _T_6_1_cf_intrVec_11 <= frontend_io_out_1_bits_cf_intrVec_11;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_brIdx <= 4'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_brIdx <= 4'h0;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_cf_brIdx <= frontend_io_out_0_bits_cf_brIdx;
            end else begin
              _T_6_1_cf_brIdx <= 4'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_cf_brIdx <= frontend_io_out_0_bits_cf_brIdx;
          end else begin
            _T_6_1_cf_brIdx <= 4'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_crossPageIPFFix <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_crossPageIPFFix <= 1'h0;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            _T_6_1_cf_crossPageIPFFix <= _T_27_cf_crossPageIPFFix;
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          _T_6_1_cf_crossPageIPFFix <= _T_27_cf_crossPageIPFFix;
        end
      end
    end
    if (reset) begin
      _T_6_1_ctrl_src1Type <= 2'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_ctrl_src1Type <= 2'h1;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_ctrl_src1Type <= frontend_io_out_0_bits_ctrl_src1Type;
            end else begin
              _T_6_1_ctrl_src1Type <= 2'h1;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_ctrl_src1Type <= frontend_io_out_0_bits_ctrl_src1Type;
          end else begin
            _T_6_1_ctrl_src1Type <= 2'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_ctrl_src2Type <= 2'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_ctrl_src2Type <= 2'h1;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_ctrl_src2Type <= frontend_io_out_0_bits_ctrl_src2Type;
            end else begin
              _T_6_1_ctrl_src2Type <= 2'h1;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_ctrl_src2Type <= frontend_io_out_0_bits_ctrl_src2Type;
          end else begin
            _T_6_1_ctrl_src2Type <= 2'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_ctrl_fuType <= 3'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_ctrl_fuType <= 3'h3;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_ctrl_fuType <= frontend_io_out_0_bits_ctrl_fuType;
            end else begin
              _T_6_1_ctrl_fuType <= 3'h3;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_ctrl_fuType <= frontend_io_out_0_bits_ctrl_fuType;
          end else begin
            _T_6_1_ctrl_fuType <= 3'h3;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_ctrl_fuOpType <= 7'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_ctrl_fuOpType <= 7'h0;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_ctrl_fuOpType <= frontend_io_out_0_bits_ctrl_fuOpType;
            end else begin
              _T_6_1_ctrl_fuOpType <= 7'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_ctrl_fuOpType <= frontend_io_out_0_bits_ctrl_fuOpType;
          end else begin
            _T_6_1_ctrl_fuOpType <= 7'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_ctrl_rfSrc1 <= 5'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_ctrl_rfSrc1 <= 5'h0;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_ctrl_rfSrc1 <= frontend_io_out_0_bits_ctrl_rfSrc1;
            end else begin
              _T_6_1_ctrl_rfSrc1 <= 5'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_ctrl_rfSrc1 <= frontend_io_out_0_bits_ctrl_rfSrc1;
          end else begin
            _T_6_1_ctrl_rfSrc1 <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_ctrl_rfSrc2 <= 5'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_ctrl_rfSrc2 <= 5'h0;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_ctrl_rfSrc2 <= frontend_io_out_0_bits_ctrl_rfSrc2;
            end else begin
              _T_6_1_ctrl_rfSrc2 <= 5'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_ctrl_rfSrc2 <= frontend_io_out_0_bits_ctrl_rfSrc2;
          end else begin
            _T_6_1_ctrl_rfSrc2 <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_ctrl_rfWen <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_ctrl_rfWen <= 1'h0;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            _T_6_1_ctrl_rfWen <= _T_27_ctrl_rfWen;
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          _T_6_1_ctrl_rfWen <= _T_27_ctrl_rfWen;
        end
      end
    end
    if (reset) begin
      _T_6_1_ctrl_rfDest <= 5'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_ctrl_rfDest <= 5'h0;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_ctrl_rfDest <= frontend_io_out_0_bits_ctrl_rfDest;
            end else begin
              _T_6_1_ctrl_rfDest <= 5'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_ctrl_rfDest <= frontend_io_out_0_bits_ctrl_rfDest;
          end else begin
            _T_6_1_ctrl_rfDest <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_ctrl_isNutCoreTrap <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_ctrl_isNutCoreTrap <= 1'h0;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            _T_6_1_ctrl_isNutCoreTrap <= _T_27_ctrl_isNutCoreTrap;
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          _T_6_1_ctrl_isNutCoreTrap <= _T_27_ctrl_isNutCoreTrap;
        end
      end
    end
    if (reset) begin
      _T_6_1_data_imm <= 64'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_data_imm <= 64'h0;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_data_imm <= frontend_io_out_0_bits_data_imm;
            end else begin
              _T_6_1_data_imm <= 64'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_data_imm <= frontend_io_out_0_bits_data_imm;
          end else begin
            _T_6_1_data_imm <= 64'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_instr <= 64'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_instr <= 64'h0;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_instr <= _T_27_cf_instr;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_instr <= _T_27_cf_instr;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_pc <= 39'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_pc <= 39'h0;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_pc <= _T_27_cf_pc;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_pc <= _T_27_cf_pc;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_pnpc <= 39'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_pnpc <= 39'h0;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_pnpc <= _T_27_cf_pnpc;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_pnpc <= _T_27_cf_pnpc;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_exceptionVec_1 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_exceptionVec_1 <= 1'h0;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_exceptionVec_1 <= _T_27_cf_exceptionVec_1;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_exceptionVec_1 <= _T_27_cf_exceptionVec_1;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_exceptionVec_2 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_exceptionVec_2 <= 1'h0;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_exceptionVec_2 <= _T_27_cf_exceptionVec_2;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_exceptionVec_2 <= _T_27_cf_exceptionVec_2;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_exceptionVec_12 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_exceptionVec_12 <= 1'h0;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_exceptionVec_12 <= _T_27_cf_exceptionVec_12;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_exceptionVec_12 <= _T_27_cf_exceptionVec_12;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_intrVec_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_intrVec_0 <= _T_6_T_29_cf_intrVec_0;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_intrVec_0 <= _T_27_cf_intrVec_0;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_intrVec_0 <= _T_27_cf_intrVec_0;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_intrVec_1 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_intrVec_1 <= _T_6_T_29_cf_intrVec_1;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_intrVec_1 <= _T_27_cf_intrVec_1;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_intrVec_1 <= _T_27_cf_intrVec_1;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_intrVec_2 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_intrVec_2 <= _T_6_T_29_cf_intrVec_2;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_intrVec_2 <= _T_27_cf_intrVec_2;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_intrVec_2 <= _T_27_cf_intrVec_2;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_intrVec_3 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_intrVec_3 <= _T_6_T_29_cf_intrVec_3;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_intrVec_3 <= _T_27_cf_intrVec_3;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_intrVec_3 <= _T_27_cf_intrVec_3;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_intrVec_4 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_intrVec_4 <= _T_6_T_29_cf_intrVec_4;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_intrVec_4 <= _T_27_cf_intrVec_4;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_intrVec_4 <= _T_27_cf_intrVec_4;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_intrVec_5 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_intrVec_5 <= _T_6_T_29_cf_intrVec_5;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_intrVec_5 <= _T_27_cf_intrVec_5;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_intrVec_5 <= _T_27_cf_intrVec_5;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_intrVec_6 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_intrVec_6 <= _T_6_T_29_cf_intrVec_6;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_intrVec_6 <= _T_27_cf_intrVec_6;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_intrVec_6 <= _T_27_cf_intrVec_6;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_intrVec_7 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_intrVec_7 <= _T_6_T_29_cf_intrVec_7;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_intrVec_7 <= _T_27_cf_intrVec_7;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_intrVec_7 <= _T_27_cf_intrVec_7;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_intrVec_8 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_intrVec_8 <= _T_6_T_29_cf_intrVec_8;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_intrVec_8 <= _T_27_cf_intrVec_8;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_intrVec_8 <= _T_27_cf_intrVec_8;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_intrVec_9 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_intrVec_9 <= _T_6_T_29_cf_intrVec_9;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_intrVec_9 <= _T_27_cf_intrVec_9;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_intrVec_9 <= _T_27_cf_intrVec_9;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_intrVec_10 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_intrVec_10 <= _T_6_T_29_cf_intrVec_10;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_intrVec_10 <= _T_27_cf_intrVec_10;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_intrVec_10 <= _T_27_cf_intrVec_10;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_intrVec_11 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_intrVec_11 <= _T_6_T_29_cf_intrVec_11;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_intrVec_11 <= _T_27_cf_intrVec_11;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_intrVec_11 <= _T_27_cf_intrVec_11;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_brIdx <= 4'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_brIdx <= 4'h0;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_brIdx <= _T_27_cf_brIdx;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_brIdx <= _T_27_cf_brIdx;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_crossPageIPFFix <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_crossPageIPFFix <= 1'h0;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_crossPageIPFFix <= _T_27_cf_crossPageIPFFix;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_crossPageIPFFix <= _T_27_cf_crossPageIPFFix;
        end
      end
    end
    if (reset) begin
      _T_6_2_ctrl_src1Type <= 2'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_ctrl_src1Type <= 2'h1;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_ctrl_src1Type <= _T_27_ctrl_src1Type;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_ctrl_src1Type <= _T_27_ctrl_src1Type;
        end
      end
    end
    if (reset) begin
      _T_6_2_ctrl_src2Type <= 2'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_ctrl_src2Type <= 2'h1;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_ctrl_src2Type <= _T_27_ctrl_src2Type;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_ctrl_src2Type <= _T_27_ctrl_src2Type;
        end
      end
    end
    if (reset) begin
      _T_6_2_ctrl_fuType <= 3'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_ctrl_fuType <= 3'h3;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_ctrl_fuType <= _T_27_ctrl_fuType;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_ctrl_fuType <= _T_27_ctrl_fuType;
        end
      end
    end
    if (reset) begin
      _T_6_2_ctrl_fuOpType <= 7'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_ctrl_fuOpType <= 7'h0;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_ctrl_fuOpType <= _T_27_ctrl_fuOpType;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_ctrl_fuOpType <= _T_27_ctrl_fuOpType;
        end
      end
    end
    if (reset) begin
      _T_6_2_ctrl_rfSrc1 <= 5'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_ctrl_rfSrc1 <= 5'h0;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_ctrl_rfSrc1 <= _T_27_ctrl_rfSrc1;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_ctrl_rfSrc1 <= _T_27_ctrl_rfSrc1;
        end
      end
    end
    if (reset) begin
      _T_6_2_ctrl_rfSrc2 <= 5'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_ctrl_rfSrc2 <= 5'h0;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_ctrl_rfSrc2 <= _T_27_ctrl_rfSrc2;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_ctrl_rfSrc2 <= _T_27_ctrl_rfSrc2;
        end
      end
    end
    if (reset) begin
      _T_6_2_ctrl_rfWen <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_ctrl_rfWen <= 1'h0;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_ctrl_rfWen <= _T_27_ctrl_rfWen;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_ctrl_rfWen <= _T_27_ctrl_rfWen;
        end
      end
    end
    if (reset) begin
      _T_6_2_ctrl_rfDest <= 5'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_ctrl_rfDest <= 5'h0;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_ctrl_rfDest <= _T_27_ctrl_rfDest;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_ctrl_rfDest <= _T_27_ctrl_rfDest;
        end
      end
    end
    if (reset) begin
      _T_6_2_ctrl_isNutCoreTrap <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_ctrl_isNutCoreTrap <= 1'h0;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_ctrl_isNutCoreTrap <= _T_27_ctrl_isNutCoreTrap;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_ctrl_isNutCoreTrap <= _T_27_ctrl_isNutCoreTrap;
        end
      end
    end
    if (reset) begin
      _T_6_2_data_imm <= 64'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_data_imm <= 64'h0;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_data_imm <= _T_27_data_imm;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_data_imm <= _T_27_data_imm;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_instr <= 64'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_instr <= 64'h0;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_instr <= _T_27_cf_instr;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_instr <= _T_27_cf_instr;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_pc <= 39'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_pc <= 39'h0;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_pc <= _T_27_cf_pc;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_pc <= _T_27_cf_pc;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_pnpc <= 39'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_pnpc <= 39'h0;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_pnpc <= _T_27_cf_pnpc;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_pnpc <= _T_27_cf_pnpc;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_exceptionVec_1 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_exceptionVec_1 <= 1'h0;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_exceptionVec_1 <= _T_27_cf_exceptionVec_1;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_exceptionVec_1 <= _T_27_cf_exceptionVec_1;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_exceptionVec_2 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_exceptionVec_2 <= 1'h0;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_exceptionVec_2 <= _T_27_cf_exceptionVec_2;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_exceptionVec_2 <= _T_27_cf_exceptionVec_2;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_exceptionVec_12 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_exceptionVec_12 <= 1'h0;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_exceptionVec_12 <= _T_27_cf_exceptionVec_12;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_exceptionVec_12 <= _T_27_cf_exceptionVec_12;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_intrVec_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_intrVec_0 <= _T_6_T_29_cf_intrVec_0;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_intrVec_0 <= _T_27_cf_intrVec_0;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_intrVec_0 <= _T_27_cf_intrVec_0;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_intrVec_1 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_intrVec_1 <= _T_6_T_29_cf_intrVec_1;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_intrVec_1 <= _T_27_cf_intrVec_1;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_intrVec_1 <= _T_27_cf_intrVec_1;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_intrVec_2 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_intrVec_2 <= _T_6_T_29_cf_intrVec_2;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_intrVec_2 <= _T_27_cf_intrVec_2;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_intrVec_2 <= _T_27_cf_intrVec_2;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_intrVec_3 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_intrVec_3 <= _T_6_T_29_cf_intrVec_3;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_intrVec_3 <= _T_27_cf_intrVec_3;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_intrVec_3 <= _T_27_cf_intrVec_3;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_intrVec_4 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_intrVec_4 <= _T_6_T_29_cf_intrVec_4;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_intrVec_4 <= _T_27_cf_intrVec_4;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_intrVec_4 <= _T_27_cf_intrVec_4;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_intrVec_5 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_intrVec_5 <= _T_6_T_29_cf_intrVec_5;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_intrVec_5 <= _T_27_cf_intrVec_5;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_intrVec_5 <= _T_27_cf_intrVec_5;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_intrVec_6 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_intrVec_6 <= _T_6_T_29_cf_intrVec_6;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_intrVec_6 <= _T_27_cf_intrVec_6;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_intrVec_6 <= _T_27_cf_intrVec_6;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_intrVec_7 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_intrVec_7 <= _T_6_T_29_cf_intrVec_7;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_intrVec_7 <= _T_27_cf_intrVec_7;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_intrVec_7 <= _T_27_cf_intrVec_7;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_intrVec_8 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_intrVec_8 <= _T_6_T_29_cf_intrVec_8;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_intrVec_8 <= _T_27_cf_intrVec_8;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_intrVec_8 <= _T_27_cf_intrVec_8;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_intrVec_9 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_intrVec_9 <= _T_6_T_29_cf_intrVec_9;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_intrVec_9 <= _T_27_cf_intrVec_9;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_intrVec_9 <= _T_27_cf_intrVec_9;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_intrVec_10 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_intrVec_10 <= _T_6_T_29_cf_intrVec_10;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_intrVec_10 <= _T_27_cf_intrVec_10;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_intrVec_10 <= _T_27_cf_intrVec_10;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_intrVec_11 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_intrVec_11 <= _T_6_T_29_cf_intrVec_11;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_intrVec_11 <= _T_27_cf_intrVec_11;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_intrVec_11 <= _T_27_cf_intrVec_11;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_brIdx <= 4'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_brIdx <= 4'h0;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_brIdx <= _T_27_cf_brIdx;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_brIdx <= _T_27_cf_brIdx;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_crossPageIPFFix <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_crossPageIPFFix <= 1'h0;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_crossPageIPFFix <= _T_27_cf_crossPageIPFFix;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_crossPageIPFFix <= _T_27_cf_crossPageIPFFix;
        end
      end
    end
    if (reset) begin
      _T_6_3_ctrl_src1Type <= 2'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_ctrl_src1Type <= 2'h1;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_ctrl_src1Type <= _T_27_ctrl_src1Type;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_ctrl_src1Type <= _T_27_ctrl_src1Type;
        end
      end
    end
    if (reset) begin
      _T_6_3_ctrl_src2Type <= 2'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_ctrl_src2Type <= 2'h1;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_ctrl_src2Type <= _T_27_ctrl_src2Type;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_ctrl_src2Type <= _T_27_ctrl_src2Type;
        end
      end
    end
    if (reset) begin
      _T_6_3_ctrl_fuType <= 3'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_ctrl_fuType <= 3'h3;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_ctrl_fuType <= _T_27_ctrl_fuType;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_ctrl_fuType <= _T_27_ctrl_fuType;
        end
      end
    end
    if (reset) begin
      _T_6_3_ctrl_fuOpType <= 7'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_ctrl_fuOpType <= 7'h0;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_ctrl_fuOpType <= _T_27_ctrl_fuOpType;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_ctrl_fuOpType <= _T_27_ctrl_fuOpType;
        end
      end
    end
    if (reset) begin
      _T_6_3_ctrl_rfSrc1 <= 5'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_ctrl_rfSrc1 <= 5'h0;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_ctrl_rfSrc1 <= _T_27_ctrl_rfSrc1;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_ctrl_rfSrc1 <= _T_27_ctrl_rfSrc1;
        end
      end
    end
    if (reset) begin
      _T_6_3_ctrl_rfSrc2 <= 5'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_ctrl_rfSrc2 <= 5'h0;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_ctrl_rfSrc2 <= _T_27_ctrl_rfSrc2;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_ctrl_rfSrc2 <= _T_27_ctrl_rfSrc2;
        end
      end
    end
    if (reset) begin
      _T_6_3_ctrl_rfWen <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_ctrl_rfWen <= 1'h0;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_ctrl_rfWen <= _T_27_ctrl_rfWen;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_ctrl_rfWen <= _T_27_ctrl_rfWen;
        end
      end
    end
    if (reset) begin
      _T_6_3_ctrl_rfDest <= 5'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_ctrl_rfDest <= 5'h0;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_ctrl_rfDest <= _T_27_ctrl_rfDest;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_ctrl_rfDest <= _T_27_ctrl_rfDest;
        end
      end
    end
    if (reset) begin
      _T_6_3_ctrl_isNutCoreTrap <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_ctrl_isNutCoreTrap <= 1'h0;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_ctrl_isNutCoreTrap <= _T_27_ctrl_isNutCoreTrap;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_ctrl_isNutCoreTrap <= _T_27_ctrl_isNutCoreTrap;
        end
      end
    end
    if (reset) begin
      _T_6_3_data_imm <= 64'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_data_imm <= 64'h0;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_data_imm <= _T_27_data_imm;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_data_imm <= _T_27_data_imm;
        end
      end
    end
    if (reset) begin
      _T_7 <= 2'h0;
    end else if (frontend_io_flushVec[1]) begin
      _T_7 <= 2'h0;
    end else if (_T_22) begin
      _T_7 <= _T_31;
    end
    if (reset) begin
      _T_8 <= 2'h0;
    end else if (frontend_io_flushVec[1]) begin
      _T_8 <= 2'h0;
    end else if (_T_44) begin
      _T_8 <= _T_46;
    end
    if (reset) begin
      _T_62 <= 64'h0;
    end else begin
      _T_62 <= _T_64;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_54) begin
          $fwrite(32'h80000002,"[DPQ] size %x head %x tail %x enq %x deq %x\n",_T_52,_T_7,_T_8,_T_19,_T_43); // @[PipelineVector.scala 77:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_54) begin
          $fwrite(32'h80000002,"[%d] NutCore: ",_T_62); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_54) begin
          $fwrite(32'h80000002,"------------------------ BACKEND ------------------------\n"); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CoherenceManager(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [3:0]  io_in_req_bits_cmd,
  input  [63:0] io_in_req_bits_wdata,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_mem_req_ready,
  output        io_out_mem_req_valid,
  output [31:0] io_out_mem_req_bits_addr,
  output [3:0]  io_out_mem_req_bits_cmd,
  output [63:0] io_out_mem_req_bits_wdata,
  output        io_out_mem_resp_ready,
  input         io_out_mem_resp_valid,
  input  [3:0]  io_out_mem_resp_bits_cmd,
  input  [63:0] io_out_mem_resp_bits_rdata,
  input         io_out_coh_req_ready,
  output        io_out_coh_req_valid,
  output [31:0] io_out_coh_req_bits_addr,
  output [63:0] io_out_coh_req_bits_wdata,
  output        io_out_coh_resp_ready,
  input         io_out_coh_resp_valid,
  input  [3:0]  io_out_coh_resp_bits_cmd,
  input  [63:0] io_out_coh_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[Coherence.scala 45:22]
  wire  inflight = state != 3'h0; // @[Coherence.scala 46:24]
  wire  _T_1 = ~io_in_req_bits_cmd[0]; // @[SimpleBus.scala 73:18]
  wire  _T_3 = ~io_in_req_bits_cmd[3]; // @[SimpleBus.scala 73:29]
  wire  _T_4 = _T_1 & _T_3; // @[SimpleBus.scala 73:26]
  wire  _T_5 = ~_T_4; // @[Coherence.scala 49:29]
  wire  _T_6 = io_in_req_valid & _T_5; // @[Coherence.scala 49:26]
  wire  _T_9 = _T_6 & _T_1; // @[Coherence.scala 49:52]
  wire  _T_10 = ~_T_9; // @[Coherence.scala 49:10]
  wire  _T_12 = _T_10 | reset; // @[Coherence.scala 49:9]
  wire  _T_13 = ~_T_12; // @[Coherence.scala 49:9]
  wire  _T_14 = ~inflight; // @[Coherence.scala 52:42]
  wire  _T_20 = _T_14 & _T_4; // @[Coherence.scala 52:52]
  reg [31:0] reqLatch_addr; // @[Reg.scala 15:16]
  reg [3:0] reqLatch_cmd; // @[Reg.scala 15:16]
  reg [63:0] reqLatch_wdata; // @[Reg.scala 15:16]
  wire  _T_23 = io_in_req_valid & _T_14; // @[Coherence.scala 65:43]
  wire  _T_25 = io_out_mem_req_ready & _T_14; // @[Coherence.scala 66:43]
  wire  _T_34 = io_out_coh_req_ready & _T_14; // @[Coherence.scala 69:43]
  wire  _GEN_5 = _T_4 & _T_23; // @[Coherence.scala 67:39]
  wire  _GEN_6 = _T_4 & _T_34; // @[Coherence.scala 67:39]
  wire  _GEN_7 = io_in_req_bits_cmd[0] & _T_23; // @[Coherence.scala 64:61]
  wire  _T_35 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_36 = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_43 = io_in_req_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_44 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_45 = io_out_coh_resp_ready & io_out_coh_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_46 = io_out_coh_resp_bits_cmd == 4'hc; // @[SimpleBus.scala 92:26]
  wire  _T_48 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_50 = io_in_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire  _T_51 = io_in_resp_valid & _T_50; // @[Coherence.scala 89:29]
  wire  _T_52 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_53 = io_out_mem_req_ready & io_out_mem_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_54 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_55 = io_out_mem_resp_ready & io_out_mem_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_56 = io_out_mem_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire  _T_57 = _T_55 & _T_56; // @[Coherence.scala 96:55]
  wire  _T_58 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire [63:0] _GEN_20 = _T_52 ? reqLatch_wdata : io_in_req_bits_wdata; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_22 = _T_52 ? reqLatch_cmd : io_in_req_bits_cmd; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_24 = _T_52 ? reqLatch_addr : io_in_req_bits_addr; // @[Conditional.scala 39:67]
  wire  _GEN_25 = _T_52 | _GEN_7; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_27 = _T_48 ? io_out_coh_resp_bits_rdata : io_out_mem_resp_bits_rdata; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_28 = _T_48 ? io_out_coh_resp_bits_cmd : io_out_mem_resp_bits_cmd; // @[Conditional.scala 39:67]
  wire  _GEN_29 = _T_48 ? io_out_coh_resp_valid : io_out_mem_resp_valid; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_32 = _T_48 ? io_in_req_bits_wdata : _GEN_20; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_34 = _T_48 ? io_in_req_bits_cmd : _GEN_22; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_36 = _T_48 ? io_in_req_bits_addr : _GEN_24; // @[Conditional.scala 39:67]
  wire  _GEN_37 = _T_48 ? _GEN_7 : _GEN_25; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_39 = _T_44 ? io_out_mem_resp_bits_rdata : _GEN_27; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_40 = _T_44 ? io_out_mem_resp_bits_cmd : _GEN_28; // @[Conditional.scala 39:67]
  wire  _GEN_41 = _T_44 ? io_out_mem_resp_valid : _GEN_29; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_43 = _T_44 ? io_in_req_bits_wdata : _GEN_32; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_45 = _T_44 ? io_in_req_bits_cmd : _GEN_34; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_47 = _T_44 ? io_in_req_bits_addr : _GEN_36; // @[Conditional.scala 39:67]
  wire  _GEN_48 = _T_44 ? _GEN_7 : _GEN_37; // @[Conditional.scala 39:67]
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _T_25 : _GEN_6; // @[Coherence.scala 62:17 Coherence.scala 66:19 Coherence.scala 69:19]
  assign io_in_resp_valid = _T_35 ? io_out_mem_resp_valid : _GEN_41; // @[Coherence.scala 72:14 Coherence.scala 88:16]
  assign io_in_resp_bits_cmd = _T_35 ? io_out_mem_resp_bits_cmd : _GEN_40; // @[Coherence.scala 72:14 Coherence.scala 88:16]
  assign io_in_resp_bits_rdata = _T_35 ? io_out_mem_resp_bits_rdata : _GEN_39; // @[Coherence.scala 72:14 Coherence.scala 88:16]
  assign io_out_mem_req_valid = _T_35 ? _GEN_7 : _GEN_48; // @[Coherence.scala 61:24 Coherence.scala 65:26 Coherence.scala 93:28]
  assign io_out_mem_req_bits_addr = _T_35 ? io_in_req_bits_addr : _GEN_47; // @[Coherence.scala 59:23 Coherence.scala 92:27]
  assign io_out_mem_req_bits_cmd = _T_35 ? io_in_req_bits_cmd : _GEN_45; // @[Coherence.scala 59:23 Coherence.scala 92:27]
  assign io_out_mem_req_bits_wdata = _T_35 ? io_in_req_bits_wdata : _GEN_43; // @[Coherence.scala 59:23 Coherence.scala 92:27]
  assign io_out_mem_resp_ready = 1'h1; // @[Coherence.scala 72:14]
  assign io_out_coh_req_valid = io_in_req_bits_cmd[0] ? 1'h0 : _GEN_5; // @[Coherence.scala 63:24 Coherence.scala 68:26]
  assign io_out_coh_req_bits_addr = io_in_req_bits_addr; // @[Coherence.scala 54:16]
  assign io_out_coh_req_bits_wdata = io_in_req_bits_wdata; // @[Coherence.scala 54:16]
  assign io_out_coh_resp_ready = 1'h1; // @[Coherence.scala 56:18 Coherence.scala 88:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  reqLatch_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reqLatch_cmd = _RAND_2[3:0];
  _RAND_3 = {2{`RANDOM}};
  reqLatch_wdata = _RAND_3[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 3'h0;
    end else if (_T_35) begin
      if (_T_36) begin
        if (_T_4) begin
          state <= 3'h1;
        end else if (_T_43) begin
          state <= 3'h5;
        end
      end
    end else if (_T_44) begin
      if (_T_45) begin
        if (_T_46) begin
          state <= 3'h2;
        end else begin
          state <= 3'h3;
        end
      end
    end else if (_T_48) begin
      if (_T_51) begin
        state <= 3'h0;
      end
    end else if (_T_52) begin
      if (_T_53) begin
        state <= 3'h4;
      end
    end else if (_T_54) begin
      if (_T_57) begin
        state <= 3'h0;
      end
    end else if (_T_58) begin
      if (_T_55) begin
        state <= 3'h0;
      end
    end
    if (_T_20) begin
      reqLatch_addr <= io_in_req_bits_addr;
    end
    if (_T_20) begin
      reqLatch_cmd <= io_in_req_bits_cmd;
    end
    if (_T_20) begin
      reqLatch_wdata <= io_in_req_bits_wdata;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Coherence.scala:49 assert(!(thisReq.valid && !thisReq.bits.isRead() && !thisReq.bits.isWrite()))\n"); // @[Coherence.scala 49:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_13) begin
          $fatal; // @[Coherence.scala 49:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module AXI42SimpleBusConverter(
  input         clock,
  input         reset,
  output        io_in_aw_ready,
  input         io_in_aw_valid,
  input  [31:0] io_in_aw_bits_addr,
  input  [7:0]  io_in_aw_bits_len,
  input  [2:0]  io_in_aw_bits_size,
  output        io_in_w_ready,
  input         io_in_w_valid,
  input  [63:0] io_in_w_bits_data,
  input  [7:0]  io_in_w_bits_strb,
  input         io_in_b_ready,
  output        io_in_b_valid,
  output        io_in_ar_ready,
  input         io_in_ar_valid,
  input  [31:0] io_in_ar_bits_addr,
  input         io_in_r_ready,
  output        io_in_r_valid,
  output [63:0] io_in_r_bits_data,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [2:0]  io_out_req_bits_size,
  output [3:0]  io_out_req_bits_cmd,
  output [7:0]  io_out_req_bits_wmask,
  output [63:0] io_out_req_bits_wdata,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [3:0]  io_out_resp_bits_cmd,
  input  [63:0] io_out_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] inflight_type; // @[ToAXI4.scala 40:30]
  wire  _T = inflight_type == 2'h0; // @[ToAXI4.scala 50:19]
  wire  _T_1 = ~_T; // @[ToAXI4.scala 53:5]
  wire  _T_2 = ~_T_1; // @[ToAXI4.scala 64:9]
  wire  _T_3 = _T_2 & io_in_ar_valid; // @[ToAXI4.scala 64:23]
  wire  _T_6 = io_out_req_ready & io_out_req_valid; // @[Decoupled.scala 40:37]
  wire [31:0] _GEN_2 = _T_3 ? io_in_ar_bits_addr : 32'h0; // @[ToAXI4.scala 64:40]
  wire [2:0] _GEN_4 = _T_3 ? 3'h2 : 3'h0; // @[ToAXI4.scala 64:40]
  wire  _T_7 = inflight_type == 2'h1; // @[ToAXI4.scala 50:19]
  wire  _T_8 = _T_7 & io_out_resp_valid; // @[ToAXI4.scala 79:27]
  wire  _T_9 = io_out_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire  _T_10 = io_in_r_ready & io_in_r_valid; // @[Decoupled.scala 40:37]
  wire  _T_12 = _T_10 & _T_9; // @[ToAXI4.scala 88:22]
  reg [31:0] aw_reg_addr; // @[ToAXI4.scala 94:19]
  reg [7:0] aw_reg_len; // @[ToAXI4.scala 94:19]
  reg [2:0] aw_reg_size; // @[ToAXI4.scala 94:19]
  reg  bresp_en; // @[ToAXI4.scala 95:25]
  wire  _T_16 = _T_2 & io_in_aw_valid; // @[ToAXI4.scala 97:23]
  wire  _T_17 = ~io_in_ar_valid; // @[ToAXI4.scala 97:42]
  wire  _T_18 = _T_16 & _T_17; // @[ToAXI4.scala 97:39]
  wire  _T_19 = io_in_aw_ready & io_in_aw_valid; // @[Decoupled.scala 40:37]
  wire  _T_20 = inflight_type == 2'h2; // @[ToAXI4.scala 50:19]
  wire  _T_21 = io_in_w_ready & io_in_w_valid; // @[Decoupled.scala 40:37]
  wire  _T_22 = _T_20 & _T_21; // @[ToAXI4.scala 105:28]
  wire  _T_23 = aw_reg_len == 8'h0; // @[ToAXI4.scala 107:31]
  wire [2:0] _T_25 = _T_23 ? 3'h1 : 3'h7; // @[ToAXI4.scala 107:19]
  wire  _GEN_37 = _T_22 | bresp_en; // @[ToAXI4.scala 105:45]
  wire  _T_26 = io_in_b_ready & io_in_b_valid; // @[Decoupled.scala 40:37]
  wire  _T_32 = _T_20 & io_in_w_valid; // @[ToAXI4.scala 127:75]
  wire  _T_38 = _T_7 & io_in_r_ready; // @[ToAXI4.scala 128:57]
  wire  _T_39 = _T_2 | _T_38; // @[ToAXI4.scala 128:35]
  wire  _T_41 = _T_20 & io_in_b_ready; // @[ToAXI4.scala 128:96]
  wire  _T_57 = io_in_ar_ready & io_in_ar_valid; // @[Decoupled.scala 40:37]
  wire  _T_62 = _T_6 & _T_2; // @[ToAXI4.scala 137:48]
  wire  _T_64 = _T_62 | reset; // @[ToAXI4.scala 137:32]
  wire  _T_65 = ~_T_64; // @[ToAXI4.scala 137:32]
  wire  _T_71 = _T_2 | reset; // @[ToAXI4.scala 138:32]
  wire  _T_72 = ~_T_71; // @[ToAXI4.scala 138:32]
  wire  _T_76 = _T_6 & _T_20; // @[ToAXI4.scala 139:48]
  wire  _T_78 = _T_76 | reset; // @[ToAXI4.scala 139:31]
  wire  _T_79 = ~_T_78; // @[ToAXI4.scala 139:31]
  wire  _T_81 = io_out_resp_ready & io_out_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_83 = _T_81 & _T_20; // @[ToAXI4.scala 140:48]
  wire  _T_85 = _T_83 | reset; // @[ToAXI4.scala 140:31]
  wire  _T_86 = ~_T_85; // @[ToAXI4.scala 140:31]
  wire  _T_90 = _T_81 & _T_7; // @[ToAXI4.scala 141:48]
  wire  _T_92 = _T_90 | reset; // @[ToAXI4.scala 141:31]
  wire  _T_93 = ~_T_92; // @[ToAXI4.scala 141:31]
  assign io_in_aw_ready = _T_2 & _T_17; // @[ToAXI4.scala 132:16]
  assign io_in_w_ready = _T_20 & io_out_req_ready; // @[ToAXI4.scala 133:16]
  assign io_in_b_valid = bresp_en & io_out_resp_valid; // @[ToAXI4.scala 134:15]
  assign io_in_ar_ready = _T_2 & io_out_req_ready; // @[ToAXI4.scala 129:16]
  assign io_in_r_valid = _T_7 & io_out_resp_valid; // @[ToAXI4.scala 80:17 ToAXI4.scala 130:15]
  assign io_in_r_bits_data = _T_8 ? io_out_resp_bits_rdata : 64'h0; // @[ToAXI4.scala 60:5 ToAXI4.scala 81:12]
  assign io_out_req_valid = _T_3 | _T_32; // @[ToAXI4.scala 65:19 ToAXI4.scala 106:19 ToAXI4.scala 127:17]
  assign io_out_req_bits_addr = _T_22 ? aw_reg_addr : _GEN_2; // @[ToAXI4.scala 59:7 ToAXI4.scala 66:14 ToAXI4.scala 109:14]
  assign io_out_req_bits_size = _T_22 ? aw_reg_size : _GEN_4; // @[ToAXI4.scala 59:7 ToAXI4.scala 69:14 ToAXI4.scala 110:14]
  assign io_out_req_bits_cmd = _T_22 ? {{1'd0}, _T_25} : 4'h0; // @[ToAXI4.scala 59:7 ToAXI4.scala 67:13 ToAXI4.scala 107:13]
  assign io_out_req_bits_wmask = _T_22 ? io_in_w_bits_strb : 8'h0; // @[ToAXI4.scala 59:7 ToAXI4.scala 71:15 ToAXI4.scala 111:15]
  assign io_out_req_bits_wdata = _T_22 ? io_in_w_bits_data : 64'h0; // @[ToAXI4.scala 59:7 ToAXI4.scala 72:15 ToAXI4.scala 112:15]
  assign io_out_resp_ready = _T_39 | _T_41; // @[ToAXI4.scala 128:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inflight_type = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  aw_reg_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  aw_reg_len = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  aw_reg_size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  bresp_en = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      inflight_type <= 2'h0;
    end else if (_T_26) begin
      inflight_type <= 2'h0;
    end else if (_T_18) begin
      if (_T_19) begin
        inflight_type <= 2'h2;
      end else if (_T_8) begin
        if (_T_12) begin
          inflight_type <= 2'h0;
        end else if (_T_3) begin
          if (_T_6) begin
            inflight_type <= 2'h1;
          end
        end
      end else if (_T_3) begin
        if (_T_6) begin
          inflight_type <= 2'h1;
        end
      end
    end else if (_T_8) begin
      if (_T_12) begin
        inflight_type <= 2'h0;
      end else if (_T_3) begin
        if (_T_6) begin
          inflight_type <= 2'h1;
        end
      end
    end else if (_T_3) begin
      if (_T_6) begin
        inflight_type <= 2'h1;
      end
    end
    if (_T_18) begin
      aw_reg_addr <= io_in_aw_bits_addr;
    end
    if (_T_18) begin
      aw_reg_len <= io_in_aw_bits_len;
    end
    if (_T_18) begin
      aw_reg_size <= io_in_aw_bits_size;
    end
    if (reset) begin
      bresp_en <= 1'h0;
    end else if (_T_26) begin
      bresp_en <= 1'h0;
    end else begin
      bresp_en <= _GEN_37;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_57 & _T_65) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:137 when (axi.ar.fire()) { assert(mem.req.fire() && !isInflight()); }\n"); // @[ToAXI4.scala 137:32]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_57 & _T_65) begin
          $fatal; // @[ToAXI4.scala 137:32]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_19 & _T_72) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:138 when (axi.aw.fire()) { assert(!isInflight()); }\n"); // @[ToAXI4.scala 138:32]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_19 & _T_72) begin
          $fatal; // @[ToAXI4.scala 138:32]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_21 & _T_79) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:139 when (axi.w.fire()) { assert(mem.req .fire() && isState(axi_write)); }\n"); // @[ToAXI4.scala 139:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_21 & _T_79) begin
          $fatal; // @[ToAXI4.scala 139:31]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_26 & _T_86) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:140 when (axi.b.fire()) { assert(mem.resp.fire() && isState(axi_write)); }\n"); // @[ToAXI4.scala 140:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_26 & _T_86) begin
          $fatal; // @[ToAXI4.scala 140:31]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & _T_93) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:141 when (axi.r.fire()) { assert(mem.resp.fire() && isState(axi_read)); }\n"); // @[ToAXI4.scala 141:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10 & _T_93) begin
          $fatal; // @[ToAXI4.scala 141:31]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Prefetcher(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [2:0]  io_in_bits_size,
  input  [3:0]  io_in_bits_cmd,
  input  [7:0]  io_in_bits_wmask,
  input  [63:0] io_in_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [2:0]  io_out_bits_size,
  output [3:0]  io_out_bits_cmd,
  output [7:0]  io_out_bits_wmask,
  output [63:0] io_out_bits_wdata,
  input         DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg  getNewReq; // @[Prefetcher.scala 37:26]
  reg [31:0] prefetchReq_addr; // @[Prefetcher.scala 38:28]
  reg [2:0] prefetchReq_size; // @[Prefetcher.scala 38:28]
  reg [7:0] prefetchReq_wmask; // @[Prefetcher.scala 38:28]
  reg [63:0] prefetchReq_wdata; // @[Prefetcher.scala 38:28]
  wire  _T_2 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  reg [31:0] lastReqAddr; // @[Reg.scala 15:16]
  wire [63:0] _GEN_9 = {{32'd0}, io_in_bits_addr}; // @[Prefetcher.scala 45:30]
  wire [63:0] _T_4 = _GEN_9 & 64'hffffffffffffffc0; // @[Prefetcher.scala 45:30]
  wire [63:0] _GEN_10 = {{32'd0}, lastReqAddr}; // @[Prefetcher.scala 45:59]
  wire [63:0] _T_5 = _GEN_10 & 64'hffffffffffffffc0; // @[Prefetcher.scala 45:59]
  wire  neqAddr = _T_4 != _T_5; // @[Prefetcher.scala 45:42]
  wire  _T_6 = ~getNewReq; // @[Prefetcher.scala 47:9]
  wire  _T_7 = ~io_in_valid; // @[Prefetcher.scala 50:20]
  wire  _T_8 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_9 = _T_7 | _T_8; // @[Prefetcher.scala 50:33]
  wire  _T_12 = _T_2 & io_in_bits_cmd[1]; // @[Prefetcher.scala 51:31]
  wire  _T_13 = _T_12 & neqAddr; // @[Prefetcher.scala 51:55]
  wire [31:0] _T_14 = prefetchReq_addr ^ 32'h30000000; // @[NutCore.scala 86:11]
  wire  _T_16 = _T_14[31:28] == 4'h0; // @[NutCore.scala 86:44]
  wire [31:0] _T_17 = prefetchReq_addr ^ 32'h40000000; // @[NutCore.scala 86:11]
  wire  _T_19 = _T_17[31:30] == 2'h0; // @[NutCore.scala 86:44]
  wire  _T_20 = _T_16 | _T_19; // @[NutCore.scala 87:15]
  wire  _T_21 = ~_T_20; // @[Prefetcher.scala 54:21]
  wire  _T_30 = _T_8 | _T_20; // @[Prefetcher.scala 56:34]
  wire  _T_31 = ~_T_30; // @[Prefetcher.scala 56:18]
  reg [63:0] _T_34; // @[GTimer.scala 24:20]
  wire [63:0] _T_36 = _T_34 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_38 = ~reset; // @[Prefetcher.scala 60:11]
  assign io_in_ready = _T_6 & _T_9; // @[Prefetcher.scala 50:17 Prefetcher.scala 55:17]
  assign io_out_valid = _T_6 ? io_in_valid : _T_21; // @[Prefetcher.scala 49:18 Prefetcher.scala 54:18]
  assign io_out_bits_addr = _T_6 ? io_in_bits_addr : prefetchReq_addr; // @[Prefetcher.scala 48:17 Prefetcher.scala 53:17]
  assign io_out_bits_size = _T_6 ? io_in_bits_size : prefetchReq_size; // @[Prefetcher.scala 48:17 Prefetcher.scala 53:17]
  assign io_out_bits_cmd = _T_6 ? io_in_bits_cmd : 4'h4; // @[Prefetcher.scala 48:17 Prefetcher.scala 53:17]
  assign io_out_bits_wmask = _T_6 ? io_in_bits_wmask : prefetchReq_wmask; // @[Prefetcher.scala 48:17 Prefetcher.scala 53:17]
  assign io_out_bits_wdata = _T_6 ? io_in_bits_wdata : prefetchReq_wdata; // @[Prefetcher.scala 48:17 Prefetcher.scala 53:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  getNewReq = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  prefetchReq_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  prefetchReq_size = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  prefetchReq_wmask = _RAND_3[7:0];
  _RAND_4 = {2{`RANDOM}};
  prefetchReq_wdata = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  lastReqAddr = _RAND_5[31:0];
  _RAND_6 = {2{`RANDOM}};
  _T_34 = _RAND_6[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      getNewReq <= 1'h0;
    end else if (_T_6) begin
      getNewReq <= _T_13;
    end else begin
      getNewReq <= _T_31;
    end
    prefetchReq_addr <= io_in_bits_addr + 32'h40;
    prefetchReq_size <= io_in_bits_size;
    prefetchReq_wmask <= io_in_bits_wmask;
    prefetchReq_wdata <= io_in_bits_wdata;
    if (_T_2) begin
      lastReqAddr <= io_in_bits_addr;
    end
    if (reset) begin
      _T_34 <= 64'h0;
    end else begin
      _T_34 <= _T_36;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_38) begin
          $fwrite(32'h80000002,"%d: [Prefetcher]: in(%d,%d), out(%d,%d), in.bits.addr = %x\n",_T_34,io_in_valid,io_in_ready,io_out_valid,io_out_ready,io_in_bits_addr); // @[Prefetcher.scala 60:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CacheStage1_2(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [2:0]  io_in_bits_size,
  input  [3:0]  io_in_bits_cmd,
  input  [7:0]  io_in_bits_wmask,
  input  [63:0] io_in_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_req_addr,
  output [2:0]  io_out_bits_req_size,
  output [3:0]  io_out_bits_req_cmd,
  output [7:0]  io_out_bits_req_wmask,
  output [63:0] io_out_bits_req_wdata,
  input         io_metaReadBus_req_ready,
  output        io_metaReadBus_req_valid,
  output [8:0]  io_metaReadBus_req_bits_setIdx,
  input  [16:0] io_metaReadBus_resp_data_0_tag,
  input         io_metaReadBus_resp_data_0_valid,
  input         io_metaReadBus_resp_data_0_dirty,
  input  [16:0] io_metaReadBus_resp_data_1_tag,
  input         io_metaReadBus_resp_data_1_valid,
  input         io_metaReadBus_resp_data_1_dirty,
  input  [16:0] io_metaReadBus_resp_data_2_tag,
  input         io_metaReadBus_resp_data_2_valid,
  input         io_metaReadBus_resp_data_2_dirty,
  input  [16:0] io_metaReadBus_resp_data_3_tag,
  input         io_metaReadBus_resp_data_3_valid,
  input         io_metaReadBus_resp_data_3_dirty,
  input         io_dataReadBus_req_ready,
  output        io_dataReadBus_req_valid,
  output [11:0] io_dataReadBus_req_bits_setIdx,
  input  [63:0] io_dataReadBus_resp_data_0_data,
  input  [63:0] io_dataReadBus_resp_data_1_data,
  input  [63:0] io_dataReadBus_resp_data_2_data,
  input  [63:0] io_dataReadBus_resp_data_3_data,
  input         DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  _T = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  reg [63:0] _T_1; // @[GTimer.scala 24:20]
  wire [63:0] _T_3 = _T_1 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_5 = _T & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  wire  _T_7 = ~reset; // @[Debug.scala 56:24]
  wire  _T_29 = io_in_valid & io_metaReadBus_req_ready; // @[Cache.scala 133:31]
  wire  _T_31 = ~io_in_valid; // @[Cache.scala 134:19]
  wire  _T_32 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_33 = _T_31 | _T_32; // @[Cache.scala 134:32]
  wire  _T_34 = _T_33 & io_metaReadBus_req_ready; // @[Cache.scala 134:50]
  reg [63:0] _T_36; // @[GTimer.scala 24:20]
  wire [63:0] _T_38 = _T_36 + 64'h1; // @[GTimer.scala 25:12]
  assign io_in_ready = _T_34 & io_dataReadBus_req_ready; // @[Cache.scala 134:15]
  assign io_out_valid = _T_29 & io_dataReadBus_req_ready; // @[Cache.scala 133:16]
  assign io_out_bits_req_addr = io_in_bits_addr; // @[Cache.scala 132:19]
  assign io_out_bits_req_size = io_in_bits_size; // @[Cache.scala 132:19]
  assign io_out_bits_req_cmd = io_in_bits_cmd; // @[Cache.scala 132:19]
  assign io_out_bits_req_wmask = io_in_bits_wmask; // @[Cache.scala 132:19]
  assign io_out_bits_req_wdata = io_in_bits_wdata; // @[Cache.scala 132:19]
  assign io_metaReadBus_req_valid = io_in_valid & io_out_ready; // @[SRAMTemplate.scala 53:20]
  assign io_metaReadBus_req_bits_setIdx = io_in_bits_addr[14:6]; // @[SRAMTemplate.scala 26:17]
  assign io_dataReadBus_req_valid = io_in_valid & io_out_ready; // @[SRAMTemplate.scala 53:20]
  assign io_dataReadBus_req_bits_setIdx = {io_in_bits_addr[14:6],io_in_bits_addr[5:3]}; // @[SRAMTemplate.scala 26:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  _T_1 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  _T_36 = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_1 <= 64'h0;
    end else begin
      _T_1 <= _T_3;
    end
    if (reset) begin
      _T_36 <= 64'h0;
    end else begin
      _T_36 <= _T_38;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5 & _T_7) begin
          $fwrite(32'h80000002,"[%d] CacheStage1_2: ",_T_1); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5 & _T_7) begin
          $fwrite(32'h80000002,"[L1$] cache stage1, addr in: %x, user: %x id: %x\n",io_in_bits_addr,1'h0,1'h0); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_7) begin
          $fwrite(32'h80000002,"[%d] CacheStage1_2: ",_T_36); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_7) begin
          $fwrite(32'h80000002,"in.ready = %d, in.valid = %d, out.valid = %d, out.ready = %d, addr = %x, cmd = %x, dataReadBus.req.valid = %d\n",io_in_ready,io_in_valid,io_out_valid,io_out_ready,io_in_bits_addr,io_in_bits_cmd,io_dataReadBus_req_valid); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CacheStage2_2(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_req_addr,
  input  [2:0]  io_in_bits_req_size,
  input  [3:0]  io_in_bits_req_cmd,
  input  [7:0]  io_in_bits_req_wmask,
  input  [63:0] io_in_bits_req_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_req_addr,
  output [2:0]  io_out_bits_req_size,
  output [3:0]  io_out_bits_req_cmd,
  output [7:0]  io_out_bits_req_wmask,
  output [63:0] io_out_bits_req_wdata,
  output [16:0] io_out_bits_metas_0_tag,
  output        io_out_bits_metas_0_valid,
  output        io_out_bits_metas_0_dirty,
  output [16:0] io_out_bits_metas_1_tag,
  output        io_out_bits_metas_1_valid,
  output        io_out_bits_metas_1_dirty,
  output [16:0] io_out_bits_metas_2_tag,
  output        io_out_bits_metas_2_valid,
  output        io_out_bits_metas_2_dirty,
  output [16:0] io_out_bits_metas_3_tag,
  output        io_out_bits_metas_3_valid,
  output        io_out_bits_metas_3_dirty,
  output [63:0] io_out_bits_datas_0_data,
  output [63:0] io_out_bits_datas_1_data,
  output [63:0] io_out_bits_datas_2_data,
  output [63:0] io_out_bits_datas_3_data,
  output        io_out_bits_hit,
  output [3:0]  io_out_bits_waymask,
  output        io_out_bits_mmio,
  output        io_out_bits_isForwardData,
  output [63:0] io_out_bits_forwardData_data_data,
  output [3:0]  io_out_bits_forwardData_waymask,
  input  [16:0] io_metaReadResp_0_tag,
  input         io_metaReadResp_0_valid,
  input         io_metaReadResp_0_dirty,
  input  [16:0] io_metaReadResp_1_tag,
  input         io_metaReadResp_1_valid,
  input         io_metaReadResp_1_dirty,
  input  [16:0] io_metaReadResp_2_tag,
  input         io_metaReadResp_2_valid,
  input         io_metaReadResp_2_dirty,
  input  [16:0] io_metaReadResp_3_tag,
  input         io_metaReadResp_3_valid,
  input         io_metaReadResp_3_dirty,
  input  [63:0] io_dataReadResp_0_data,
  input  [63:0] io_dataReadResp_1_data,
  input  [63:0] io_dataReadResp_2_data,
  input  [63:0] io_dataReadResp_3_data,
  input         io_metaWriteBus_req_valid,
  input  [8:0]  io_metaWriteBus_req_bits_setIdx,
  input  [16:0] io_metaWriteBus_req_bits_data_tag,
  input         io_metaWriteBus_req_bits_data_dirty,
  input  [3:0]  io_metaWriteBus_req_bits_waymask,
  input         io_dataWriteBus_req_valid,
  input  [11:0] io_dataWriteBus_req_bits_setIdx,
  input  [63:0] io_dataWriteBus_req_bits_data_data,
  input  [3:0]  io_dataWriteBus_req_bits_waymask,
  input         DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[Cache.scala 162:31]
  wire [8:0] addr_index = io_in_bits_req_addr[14:6]; // @[Cache.scala 162:31]
  wire [16:0] addr_tag = io_in_bits_req_addr[31:15]; // @[Cache.scala 162:31]
  wire  _T_5 = io_in_valid & io_metaWriteBus_req_valid; // @[Cache.scala 164:35]
  wire  _T_12 = io_metaWriteBus_req_bits_setIdx == addr_index; // @[Cache.scala 164:99]
  wire  isForwardMeta = _T_5 & _T_12; // @[Cache.scala 164:64]
  reg  isForwardMetaReg; // @[Cache.scala 165:33]
  wire  _GEN_0 = isForwardMeta | isForwardMetaReg; // @[Cache.scala 166:24]
  wire  _T_13 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire  _T_14 = ~io_in_valid; // @[Cache.scala 167:25]
  wire  _T_15 = _T_13 | _T_14; // @[Cache.scala 167:22]
  reg [16:0] forwardMetaReg_data_tag; // @[Reg.scala 15:16]
  reg  forwardMetaReg_data_dirty; // @[Reg.scala 15:16]
  reg [3:0] forwardMetaReg_waymask; // @[Reg.scala 15:16]
  wire [3:0] _GEN_2 = isForwardMeta ? io_metaWriteBus_req_bits_waymask : forwardMetaReg_waymask; // @[Reg.scala 16:19]
  wire  _GEN_3 = isForwardMeta ? io_metaWriteBus_req_bits_data_dirty : forwardMetaReg_data_dirty; // @[Reg.scala 16:19]
  wire [16:0] _GEN_5 = isForwardMeta ? io_metaWriteBus_req_bits_data_tag : forwardMetaReg_data_tag; // @[Reg.scala 16:19]
  wire  pickForwardMeta = isForwardMetaReg | isForwardMeta; // @[Cache.scala 171:42]
  wire  forwardWaymask_0 = _GEN_2[0]; // @[Cache.scala 173:61]
  wire  forwardWaymask_1 = _GEN_2[1]; // @[Cache.scala 173:61]
  wire  forwardWaymask_2 = _GEN_2[2]; // @[Cache.scala 173:61]
  wire  forwardWaymask_3 = _GEN_2[3]; // @[Cache.scala 173:61]
  wire  _T_16 = pickForwardMeta & forwardWaymask_0; // @[Cache.scala 175:39]
  wire [16:0] metaWay_0_tag = _T_16 ? _GEN_5 : io_metaReadResp_0_tag; // @[Cache.scala 175:22]
  wire  metaWay_0_valid = _T_16 | io_metaReadResp_0_valid; // @[Cache.scala 175:22]
  wire  _T_18 = pickForwardMeta & forwardWaymask_1; // @[Cache.scala 175:39]
  wire [16:0] metaWay_1_tag = _T_18 ? _GEN_5 : io_metaReadResp_1_tag; // @[Cache.scala 175:22]
  wire  metaWay_1_valid = _T_18 | io_metaReadResp_1_valid; // @[Cache.scala 175:22]
  wire  _T_20 = pickForwardMeta & forwardWaymask_2; // @[Cache.scala 175:39]
  wire [16:0] metaWay_2_tag = _T_20 ? _GEN_5 : io_metaReadResp_2_tag; // @[Cache.scala 175:22]
  wire  metaWay_2_valid = _T_20 | io_metaReadResp_2_valid; // @[Cache.scala 175:22]
  wire  _T_22 = pickForwardMeta & forwardWaymask_3; // @[Cache.scala 175:39]
  wire [16:0] metaWay_3_tag = _T_22 ? _GEN_5 : io_metaReadResp_3_tag; // @[Cache.scala 175:22]
  wire  metaWay_3_valid = _T_22 | io_metaReadResp_3_valid; // @[Cache.scala 175:22]
  wire  _T_24 = metaWay_0_tag == addr_tag; // @[Cache.scala 178:59]
  wire  _T_25 = metaWay_0_valid & _T_24; // @[Cache.scala 178:49]
  wire  _T_26 = _T_25 & io_in_valid; // @[Cache.scala 178:73]
  wire  _T_27 = metaWay_1_tag == addr_tag; // @[Cache.scala 178:59]
  wire  _T_28 = metaWay_1_valid & _T_27; // @[Cache.scala 178:49]
  wire  _T_29 = _T_28 & io_in_valid; // @[Cache.scala 178:73]
  wire  _T_30 = metaWay_2_tag == addr_tag; // @[Cache.scala 178:59]
  wire  _T_31 = metaWay_2_valid & _T_30; // @[Cache.scala 178:49]
  wire  _T_32 = _T_31 & io_in_valid; // @[Cache.scala 178:73]
  wire  _T_33 = metaWay_3_tag == addr_tag; // @[Cache.scala 178:59]
  wire  _T_34 = metaWay_3_valid & _T_33; // @[Cache.scala 178:49]
  wire  _T_35 = _T_34 & io_in_valid; // @[Cache.scala 178:73]
  wire [3:0] hitVec = {_T_35,_T_32,_T_29,_T_26}; // @[Cache.scala 178:90]
  reg [63:0] _T_39; // @[LFSR64.scala 25:23]
  wire  _T_42 = _T_39[0] ^ _T_39[1]; // @[LFSR64.scala 26:23]
  wire  _T_44 = _T_42 ^ _T_39[3]; // @[LFSR64.scala 26:33]
  wire  _T_46 = _T_44 ^ _T_39[4]; // @[LFSR64.scala 26:43]
  wire  _T_47 = _T_39 == 64'h0; // @[LFSR64.scala 28:24]
  wire [63:0] _T_49 = {_T_46,_T_39[63:1]}; // @[Cat.scala 29:58]
  wire [3:0] victimWaymask = 4'h1 << _T_39[1:0]; // @[Cache.scala 179:42]
  wire  _T_52 = ~metaWay_0_valid; // @[Cache.scala 181:45]
  wire  _T_53 = ~metaWay_1_valid; // @[Cache.scala 181:45]
  wire  _T_54 = ~metaWay_2_valid; // @[Cache.scala 181:45]
  wire  _T_55 = ~metaWay_3_valid; // @[Cache.scala 181:45]
  wire [3:0] invalidVec = {_T_55,_T_54,_T_53,_T_52}; // @[Cache.scala 181:56]
  wire  hasInvalidWay = |invalidVec; // @[Cache.scala 182:34]
  wire  _T_59 = invalidVec >= 4'h8; // @[Cache.scala 183:45]
  wire  _T_60 = invalidVec >= 4'h4; // @[Cache.scala 184:20]
  wire  _T_61 = invalidVec >= 4'h2; // @[Cache.scala 185:20]
  wire [1:0] _T_62 = _T_61 ? 2'h2 : 2'h1; // @[Cache.scala 185:8]
  wire [2:0] _T_63 = _T_60 ? 3'h4 : {{1'd0}, _T_62}; // @[Cache.scala 184:8]
  wire [3:0] refillInvalidWaymask = _T_59 ? 4'h8 : {{1'd0}, _T_63}; // @[Cache.scala 183:33]
  wire [3:0] _T_64 = hasInvalidWay ? refillInvalidWaymask : victimWaymask; // @[Cache.scala 188:49]
  wire [3:0] waymask = io_out_bits_hit ? hitVec : _T_64; // @[Cache.scala 188:20]
  wire [1:0] _T_69 = waymask[0] + waymask[1]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_71 = waymask[2] + waymask[3]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_73 = _T_69 + _T_71; // @[Bitwise.scala 47:55]
  wire  _T_75 = _T_73 > 3'h1; // @[Cache.scala 189:26]
  reg [63:0] _T_76; // @[GTimer.scala 24:20]
  wire [63:0] _T_78 = _T_76 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_82 = ~reset; // @[Debug.scala 56:24]
  reg [63:0] _T_85; // @[GTimer.scala 24:20]
  wire [63:0] _T_87 = _T_85 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_94; // @[GTimer.scala 24:20]
  wire [63:0] _T_96 = _T_94 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_103; // @[GTimer.scala 24:20]
  wire [63:0] _T_105 = _T_103 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_112; // @[GTimer.scala 24:20]
  wire [63:0] _T_114 = _T_112 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_121; // @[GTimer.scala 24:20]
  wire [63:0] _T_123 = _T_121 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_130; // @[GTimer.scala 24:20]
  wire [63:0] _T_132 = _T_130 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_139; // @[GTimer.scala 24:20]
  wire [63:0] _T_141 = _T_139 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_148; // @[GTimer.scala 24:20]
  wire [63:0] _T_150 = _T_148 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_157; // @[GTimer.scala 24:20]
  wire [63:0] _T_159 = _T_157 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_177; // @[GTimer.scala 24:20]
  wire [63:0] _T_179 = _T_177 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_197 = io_in_valid & _T_75; // @[Cache.scala 196:24]
  wire  _T_198 = ~_T_197; // @[Cache.scala 196:10]
  wire  _T_200 = _T_198 | reset; // @[Cache.scala 196:9]
  wire  _T_201 = ~_T_200; // @[Cache.scala 196:9]
  wire  _T_202 = |hitVec; // @[Cache.scala 199:44]
  wire [31:0] _T_204 = io_in_bits_req_addr ^ 32'h30000000; // @[NutCore.scala 86:11]
  wire  _T_206 = _T_204[31:28] == 4'h0; // @[NutCore.scala 86:44]
  wire [31:0] _T_207 = io_in_bits_req_addr ^ 32'h40000000; // @[NutCore.scala 86:11]
  wire  _T_209 = _T_207[31:30] == 2'h0; // @[NutCore.scala 86:44]
  wire [11:0] _T_223 = {addr_index,addr_wordIndex}; // @[Cat.scala 29:58]
  wire  _T_224 = io_dataWriteBus_req_bits_setIdx == _T_223; // @[Cache.scala 205:30]
  wire  _T_225 = io_dataWriteBus_req_valid & _T_224; // @[Cache.scala 205:13]
  wire  isForwardData = io_in_valid & _T_225; // @[Cache.scala 204:35]
  reg  isForwardDataReg; // @[Cache.scala 207:33]
  wire  _GEN_8 = isForwardData | isForwardDataReg; // @[Cache.scala 208:24]
  reg [63:0] forwardDataReg_data_data; // @[Reg.scala 15:16]
  reg [3:0] forwardDataReg_waymask; // @[Reg.scala 15:16]
  wire  _T_232 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  reg [63:0] _T_235; // @[GTimer.scala 24:20]
  wire [63:0] _T_237 = _T_235 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_250; // @[GTimer.scala 24:20]
  wire [63:0] _T_252 = _T_250 + 64'h1; // @[GTimer.scala 25:12]
  wire  _GEN_13 = _T_75 & DISPLAY_ENABLE; // @[Debug.scala 56:24]
  assign io_in_ready = _T_14 | _T_232; // @[Cache.scala 216:15]
  assign io_out_valid = io_in_valid; // @[Cache.scala 215:16]
  assign io_out_bits_req_addr = io_in_bits_req_addr; // @[Cache.scala 214:19]
  assign io_out_bits_req_size = io_in_bits_req_size; // @[Cache.scala 214:19]
  assign io_out_bits_req_cmd = io_in_bits_req_cmd; // @[Cache.scala 214:19]
  assign io_out_bits_req_wmask = io_in_bits_req_wmask; // @[Cache.scala 214:19]
  assign io_out_bits_req_wdata = io_in_bits_req_wdata; // @[Cache.scala 214:19]
  assign io_out_bits_metas_0_tag = _T_16 ? _GEN_5 : io_metaReadResp_0_tag; // @[Cache.scala 198:21]
  assign io_out_bits_metas_0_valid = _T_16 | io_metaReadResp_0_valid; // @[Cache.scala 198:21]
  assign io_out_bits_metas_0_dirty = _T_16 ? _GEN_3 : io_metaReadResp_0_dirty; // @[Cache.scala 198:21]
  assign io_out_bits_metas_1_tag = _T_18 ? _GEN_5 : io_metaReadResp_1_tag; // @[Cache.scala 198:21]
  assign io_out_bits_metas_1_valid = _T_18 | io_metaReadResp_1_valid; // @[Cache.scala 198:21]
  assign io_out_bits_metas_1_dirty = _T_18 ? _GEN_3 : io_metaReadResp_1_dirty; // @[Cache.scala 198:21]
  assign io_out_bits_metas_2_tag = _T_20 ? _GEN_5 : io_metaReadResp_2_tag; // @[Cache.scala 198:21]
  assign io_out_bits_metas_2_valid = _T_20 | io_metaReadResp_2_valid; // @[Cache.scala 198:21]
  assign io_out_bits_metas_2_dirty = _T_20 ? _GEN_3 : io_metaReadResp_2_dirty; // @[Cache.scala 198:21]
  assign io_out_bits_metas_3_tag = _T_22 ? _GEN_5 : io_metaReadResp_3_tag; // @[Cache.scala 198:21]
  assign io_out_bits_metas_3_valid = _T_22 | io_metaReadResp_3_valid; // @[Cache.scala 198:21]
  assign io_out_bits_metas_3_dirty = _T_22 ? _GEN_3 : io_metaReadResp_3_dirty; // @[Cache.scala 198:21]
  assign io_out_bits_datas_0_data = io_dataReadResp_0_data; // @[Cache.scala 201:21]
  assign io_out_bits_datas_1_data = io_dataReadResp_1_data; // @[Cache.scala 201:21]
  assign io_out_bits_datas_2_data = io_dataReadResp_2_data; // @[Cache.scala 201:21]
  assign io_out_bits_datas_3_data = io_dataReadResp_3_data; // @[Cache.scala 201:21]
  assign io_out_bits_hit = io_in_valid & _T_202; // @[Cache.scala 199:19]
  assign io_out_bits_waymask = io_out_bits_hit ? hitVec : _T_64; // @[Cache.scala 200:23]
  assign io_out_bits_mmio = _T_206 | _T_209; // @[Cache.scala 202:20]
  assign io_out_bits_isForwardData = isForwardDataReg | isForwardData; // @[Cache.scala 211:29]
  assign io_out_bits_forwardData_data_data = isForwardData ? io_dataWriteBus_req_bits_data_data : forwardDataReg_data_data; // @[Cache.scala 212:27]
  assign io_out_bits_forwardData_waymask = isForwardData ? io_dataWriteBus_req_bits_waymask : forwardDataReg_waymask; // @[Cache.scala 212:27]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  isForwardMetaReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  forwardMetaReg_data_tag = _RAND_1[16:0];
  _RAND_2 = {1{`RANDOM}};
  forwardMetaReg_data_dirty = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  forwardMetaReg_waymask = _RAND_3[3:0];
  _RAND_4 = {2{`RANDOM}};
  _T_39 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  _T_76 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  _T_85 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  _T_94 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  _T_103 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  _T_112 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  _T_121 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  _T_130 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  _T_139 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  _T_148 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  _T_157 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  _T_177 = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  isForwardDataReg = _RAND_16[0:0];
  _RAND_17 = {2{`RANDOM}};
  forwardDataReg_data_data = _RAND_17[63:0];
  _RAND_18 = {1{`RANDOM}};
  forwardDataReg_waymask = _RAND_18[3:0];
  _RAND_19 = {2{`RANDOM}};
  _T_235 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  _T_250 = _RAND_20[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      isForwardMetaReg <= 1'h0;
    end else if (_T_15) begin
      isForwardMetaReg <= 1'h0;
    end else begin
      isForwardMetaReg <= _GEN_0;
    end
    if (isForwardMeta) begin
      forwardMetaReg_data_tag <= io_metaWriteBus_req_bits_data_tag;
    end
    if (isForwardMeta) begin
      forwardMetaReg_data_dirty <= io_metaWriteBus_req_bits_data_dirty;
    end
    if (isForwardMeta) begin
      forwardMetaReg_waymask <= io_metaWriteBus_req_bits_waymask;
    end
    if (reset) begin
      _T_39 <= 64'h1234567887654321;
    end else if (_T_47) begin
      _T_39 <= 64'h1;
    end else begin
      _T_39 <= _T_49;
    end
    if (reset) begin
      _T_76 <= 64'h0;
    end else begin
      _T_76 <= _T_78;
    end
    if (reset) begin
      _T_85 <= 64'h0;
    end else begin
      _T_85 <= _T_87;
    end
    if (reset) begin
      _T_94 <= 64'h0;
    end else begin
      _T_94 <= _T_96;
    end
    if (reset) begin
      _T_103 <= 64'h0;
    end else begin
      _T_103 <= _T_105;
    end
    if (reset) begin
      _T_112 <= 64'h0;
    end else begin
      _T_112 <= _T_114;
    end
    if (reset) begin
      _T_121 <= 64'h0;
    end else begin
      _T_121 <= _T_123;
    end
    if (reset) begin
      _T_130 <= 64'h0;
    end else begin
      _T_130 <= _T_132;
    end
    if (reset) begin
      _T_139 <= 64'h0;
    end else begin
      _T_139 <= _T_141;
    end
    if (reset) begin
      _T_148 <= 64'h0;
    end else begin
      _T_148 <= _T_150;
    end
    if (reset) begin
      _T_157 <= 64'h0;
    end else begin
      _T_157 <= _T_159;
    end
    if (reset) begin
      _T_177 <= 64'h0;
    end else begin
      _T_177 <= _T_179;
    end
    if (reset) begin
      isForwardDataReg <= 1'h0;
    end else if (_T_15) begin
      isForwardDataReg <= 1'h0;
    end else begin
      isForwardDataReg <= _GEN_8;
    end
    if (isForwardData) begin
      forwardDataReg_data_data <= io_dataWriteBus_req_bits_data_data;
    end
    if (isForwardData) begin
      forwardDataReg_waymask <= io_dataWriteBus_req_bits_waymask;
    end
    if (reset) begin
      _T_235 <= 64'h0;
    end else begin
      _T_235 <= _T_237;
    end
    if (reset) begin
      _T_250 <= 64'h0;
    end else begin
      _T_250 <= _T_252;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_2: ",_T_76); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] metaWay %x metat %x reqt %x\n",metaWay_0_valid,metaWay_0_tag,addr_tag); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_2: ",_T_85); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] metaWay %x metat %x reqt %x\n",metaWay_1_valid,metaWay_1_tag,addr_tag); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_2: ",_T_94); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] metaWay %x metat %x reqt %x\n",metaWay_2_valid,metaWay_2_tag,addr_tag); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_2: ",_T_103); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] metaWay %x metat %x reqt %x\n",metaWay_3_valid,metaWay_3_tag,addr_tag); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_2: ",_T_112); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] metaReadResp %x metat %x reqt %x\n",io_metaReadResp_0_valid,io_metaReadResp_0_tag,addr_tag); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_2: ",_T_121); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] metaReadResp %x metat %x reqt %x\n",io_metaReadResp_1_valid,io_metaReadResp_1_tag,addr_tag); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_2: ",_T_130); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] metaReadResp %x metat %x reqt %x\n",io_metaReadResp_2_valid,io_metaReadResp_2_tag,addr_tag); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_2: ",_T_139); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] metaReadResp %x metat %x reqt %x\n",io_metaReadResp_3_valid,io_metaReadResp_3_tag,addr_tag); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_2: ",_T_148); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] forwardMetaReg isForwardMetaReg %x %x metat %x wm %b\n",isForwardMetaReg,1'h1,forwardMetaReg_data_tag,forwardMetaReg_waymask); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_2: ",_T_157); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] forwardMeta isForwardMeta %x %x metat %x wm %b\n",isForwardMeta,1'h1,io_metaWriteBus_req_bits_data_tag,io_metaWriteBus_req_bits_waymask); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_2: ",_T_177); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_13 & _T_82) begin
          $fwrite(32'h80000002,"[ERROR] hit %b wmask %b hitvec %b\n",io_out_bits_hit,_GEN_2,hitVec); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_201) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Cache.scala:196 assert(!(io.in.valid && PopCount(waymask) > 1.U))\n"); // @[Cache.scala 196:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_201) begin
          $fatal; // @[Cache.scala 196:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_2: ",_T_235); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_82) begin
          $fwrite(32'h80000002,"[isFD:%d isFDreg:%d inFire:%d invalid:%d \n",isForwardData,isForwardDataReg,_T_13,io_in_valid); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_82) begin
          $fwrite(32'h80000002,"[%d] CacheStage2_2: ",_T_250); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_82) begin
          $fwrite(32'h80000002,"[isFM:%d isFMreg:%d metawreq:%x widx:%x ridx:%x \n",isForwardMeta,isForwardMetaReg,io_metaWriteBus_req_valid,io_metaWriteBus_req_bits_setIdx,addr_index); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Arbiter_10(
  input         io_in_0_valid,
  input  [8:0]  io_in_0_bits_setIdx,
  input  [16:0] io_in_0_bits_data_tag,
  input  [3:0]  io_in_0_bits_waymask,
  input         io_in_1_valid,
  input  [8:0]  io_in_1_bits_setIdx,
  input  [16:0] io_in_1_bits_data_tag,
  input         io_in_1_bits_data_dirty,
  input  [3:0]  io_in_1_bits_waymask,
  output        io_out_valid,
  output [8:0]  io_out_bits_setIdx,
  output [16:0] io_out_bits_data_tag,
  output        io_out_bits_data_dirty,
  output [3:0]  io_out_bits_waymask
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  wire  _T_2 = ~grant_1; // @[Arbiter.scala 135:19]
  assign io_out_valid = _T_2 | io_in_1_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_data_tag = io_in_0_valid ? io_in_0_bits_data_tag : io_in_1_bits_data_tag; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_data_dirty = io_in_0_valid | io_in_1_bits_data_dirty; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_waymask = io_in_0_valid ? io_in_0_bits_waymask : io_in_1_bits_waymask; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
endmodule
module Arbiter_11(
  input         io_in_0_valid,
  input  [11:0] io_in_0_bits_setIdx,
  input  [63:0] io_in_0_bits_data_data,
  input  [3:0]  io_in_0_bits_waymask,
  input         io_in_1_valid,
  input  [11:0] io_in_1_bits_setIdx,
  input  [63:0] io_in_1_bits_data_data,
  input  [3:0]  io_in_1_bits_waymask,
  output        io_out_valid,
  output [11:0] io_out_bits_setIdx,
  output [63:0] io_out_bits_data_data,
  output [3:0]  io_out_bits_waymask
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  wire  _T_2 = ~grant_1; // @[Arbiter.scala 135:19]
  assign io_out_valid = _T_2 | io_in_1_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_data_data = io_in_0_valid ? io_in_0_bits_data_data : io_in_1_bits_data_data; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_waymask = io_in_0_valid ? io_in_0_bits_waymask : io_in_1_bits_waymask; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
endmodule
module CacheStage3_2(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_req_addr,
  input  [2:0]  io_in_bits_req_size,
  input  [3:0]  io_in_bits_req_cmd,
  input  [7:0]  io_in_bits_req_wmask,
  input  [63:0] io_in_bits_req_wdata,
  input  [16:0] io_in_bits_metas_0_tag,
  input         io_in_bits_metas_0_valid,
  input         io_in_bits_metas_0_dirty,
  input  [16:0] io_in_bits_metas_1_tag,
  input         io_in_bits_metas_1_valid,
  input         io_in_bits_metas_1_dirty,
  input  [16:0] io_in_bits_metas_2_tag,
  input         io_in_bits_metas_2_valid,
  input         io_in_bits_metas_2_dirty,
  input  [16:0] io_in_bits_metas_3_tag,
  input         io_in_bits_metas_3_valid,
  input         io_in_bits_metas_3_dirty,
  input  [63:0] io_in_bits_datas_0_data,
  input  [63:0] io_in_bits_datas_1_data,
  input  [63:0] io_in_bits_datas_2_data,
  input  [63:0] io_in_bits_datas_3_data,
  input         io_in_bits_hit,
  input  [3:0]  io_in_bits_waymask,
  input         io_in_bits_mmio,
  input         io_in_bits_isForwardData,
  input  [63:0] io_in_bits_forwardData_data_data,
  input  [3:0]  io_in_bits_forwardData_waymask,
  input         io_out_ready,
  output        io_out_valid,
  output [3:0]  io_out_bits_cmd,
  output [63:0] io_out_bits_rdata,
  output        io_isFinish,
  input         io_dataReadBus_req_ready,
  output        io_dataReadBus_req_valid,
  output [11:0] io_dataReadBus_req_bits_setIdx,
  input  [63:0] io_dataReadBus_resp_data_0_data,
  input  [63:0] io_dataReadBus_resp_data_1_data,
  input  [63:0] io_dataReadBus_resp_data_2_data,
  input  [63:0] io_dataReadBus_resp_data_3_data,
  output        io_dataWriteBus_req_valid,
  output [11:0] io_dataWriteBus_req_bits_setIdx,
  output [63:0] io_dataWriteBus_req_bits_data_data,
  output [3:0]  io_dataWriteBus_req_bits_waymask,
  output        io_metaWriteBus_req_valid,
  output [8:0]  io_metaWriteBus_req_bits_setIdx,
  output [16:0] io_metaWriteBus_req_bits_data_tag,
  output        io_metaWriteBus_req_bits_data_valid,
  output        io_metaWriteBus_req_bits_data_dirty,
  output [3:0]  io_metaWriteBus_req_bits_waymask,
  input         io_mem_req_ready,
  output        io_mem_req_valid,
  output [31:0] io_mem_req_bits_addr,
  output [2:0]  io_mem_req_bits_size,
  output [3:0]  io_mem_req_bits_cmd,
  output [7:0]  io_mem_req_bits_wmask,
  output [63:0] io_mem_req_bits_wdata,
  output        io_mem_resp_ready,
  input         io_mem_resp_valid,
  input  [3:0]  io_mem_resp_bits_cmd,
  input  [63:0] io_mem_resp_bits_rdata,
  output        io_cohResp_valid,
  output        io_dataReadRespToL1,
  input         DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
`endif // RANDOMIZE_REG_INIT
  wire  metaWriteArb_io_in_0_valid; // @[Cache.scala 241:28]
  wire [8:0] metaWriteArb_io_in_0_bits_setIdx; // @[Cache.scala 241:28]
  wire [16:0] metaWriteArb_io_in_0_bits_data_tag; // @[Cache.scala 241:28]
  wire [3:0] metaWriteArb_io_in_0_bits_waymask; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_in_1_valid; // @[Cache.scala 241:28]
  wire [8:0] metaWriteArb_io_in_1_bits_setIdx; // @[Cache.scala 241:28]
  wire [16:0] metaWriteArb_io_in_1_bits_data_tag; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_in_1_bits_data_dirty; // @[Cache.scala 241:28]
  wire [3:0] metaWriteArb_io_in_1_bits_waymask; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_out_valid; // @[Cache.scala 241:28]
  wire [8:0] metaWriteArb_io_out_bits_setIdx; // @[Cache.scala 241:28]
  wire [16:0] metaWriteArb_io_out_bits_data_tag; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_out_bits_data_dirty; // @[Cache.scala 241:28]
  wire [3:0] metaWriteArb_io_out_bits_waymask; // @[Cache.scala 241:28]
  wire  dataWriteArb_io_in_0_valid; // @[Cache.scala 242:28]
  wire [11:0] dataWriteArb_io_in_0_bits_setIdx; // @[Cache.scala 242:28]
  wire [63:0] dataWriteArb_io_in_0_bits_data_data; // @[Cache.scala 242:28]
  wire [3:0] dataWriteArb_io_in_0_bits_waymask; // @[Cache.scala 242:28]
  wire  dataWriteArb_io_in_1_valid; // @[Cache.scala 242:28]
  wire [11:0] dataWriteArb_io_in_1_bits_setIdx; // @[Cache.scala 242:28]
  wire [63:0] dataWriteArb_io_in_1_bits_data_data; // @[Cache.scala 242:28]
  wire [3:0] dataWriteArb_io_in_1_bits_waymask; // @[Cache.scala 242:28]
  wire  dataWriteArb_io_out_valid; // @[Cache.scala 242:28]
  wire [11:0] dataWriteArb_io_out_bits_setIdx; // @[Cache.scala 242:28]
  wire [63:0] dataWriteArb_io_out_bits_data_data; // @[Cache.scala 242:28]
  wire [3:0] dataWriteArb_io_out_bits_waymask; // @[Cache.scala 242:28]
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[Cache.scala 245:31]
  wire [8:0] addr_index = io_in_bits_req_addr[14:6]; // @[Cache.scala 245:31]
  wire [16:0] addr_tag = io_in_bits_req_addr[31:15]; // @[Cache.scala 245:31]
  wire  mmio = io_in_valid & io_in_bits_mmio; // @[Cache.scala 246:26]
  wire  hit = io_in_valid & io_in_bits_hit; // @[Cache.scala 247:25]
  wire  _T_5 = ~io_in_bits_hit; // @[Cache.scala 248:29]
  wire  miss = io_in_valid & _T_5; // @[Cache.scala 248:26]
  wire  _T_7 = io_in_bits_req_cmd == 4'h8; // @[SimpleBus.scala 79:23]
  wire  probe = io_in_valid & _T_7; // @[Cache.scala 249:39]
  wire  _T_8 = io_in_bits_req_cmd == 4'h2; // @[SimpleBus.scala 76:27]
  wire  hitReadBurst = hit & _T_8; // @[Cache.scala 250:26]
  wire [18:0] _T_14 = {io_in_bits_metas_0_tag,io_in_bits_metas_0_valid,io_in_bits_metas_0_dirty}; // @[Mux.scala 27:72]
  wire [18:0] _T_15 = io_in_bits_waymask[0] ? _T_14 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_17 = {io_in_bits_metas_1_tag,io_in_bits_metas_1_valid,io_in_bits_metas_1_dirty}; // @[Mux.scala 27:72]
  wire [18:0] _T_18 = io_in_bits_waymask[1] ? _T_17 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_20 = {io_in_bits_metas_2_tag,io_in_bits_metas_2_valid,io_in_bits_metas_2_dirty}; // @[Mux.scala 27:72]
  wire [18:0] _T_21 = io_in_bits_waymask[2] ? _T_20 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_23 = {io_in_bits_metas_3_tag,io_in_bits_metas_3_valid,io_in_bits_metas_3_dirty}; // @[Mux.scala 27:72]
  wire [18:0] _T_24 = io_in_bits_waymask[3] ? _T_23 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_25 = _T_15 | _T_18; // @[Mux.scala 27:72]
  wire [18:0] _T_26 = _T_25 | _T_21; // @[Mux.scala 27:72]
  wire [18:0] _T_27 = _T_26 | _T_24; // @[Mux.scala 27:72]
  wire  meta_dirty = _T_27[0]; // @[Mux.scala 27:72]
  wire [16:0] meta_tag = _T_27[18:2]; // @[Mux.scala 27:72]
  wire  _T_32 = mmio & hit; // @[Cache.scala 252:17]
  wire  _T_33 = ~_T_32; // @[Cache.scala 252:10]
  wire  _T_35 = _T_33 | reset; // @[Cache.scala 252:9]
  wire  _T_36 = ~_T_35; // @[Cache.scala 252:9]
  wire  _T_37 = io_in_bits_waymask == io_in_bits_forwardData_waymask; // @[Cache.scala 260:71]
  wire  useForwardData = io_in_bits_isForwardData & _T_37; // @[Cache.scala 260:49]
  wire [63:0] _T_42 = io_in_bits_waymask[0] ? io_in_bits_datas_0_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_43 = io_in_bits_waymask[1] ? io_in_bits_datas_1_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_44 = io_in_bits_waymask[2] ? io_in_bits_datas_2_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_45 = io_in_bits_waymask[3] ? io_in_bits_datas_3_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_46 = _T_42 | _T_43; // @[Mux.scala 27:72]
  wire [63:0] _T_47 = _T_46 | _T_44; // @[Mux.scala 27:72]
  wire [63:0] _T_48 = _T_47 | _T_45; // @[Mux.scala 27:72]
  wire [63:0] dataRead = useForwardData ? io_in_bits_forwardData_data_data : _T_48; // @[Cache.scala 262:21]
  wire [7:0] _T_64 = io_in_bits_req_wmask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_66 = io_in_bits_req_wmask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_68 = io_in_bits_req_wmask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_70 = io_in_bits_req_wmask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_72 = io_in_bits_req_wmask[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_74 = io_in_bits_req_wmask[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_76 = io_in_bits_req_wmask[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_78 = io_in_bits_req_wmask[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_85 = {_T_78,_T_76,_T_74,_T_72,_T_70,_T_68,_T_66,_T_64}; // @[Cat.scala 29:58]
  wire [63:0] wordMask = io_in_bits_req_cmd[0] ? _T_85 : 64'h0; // @[Cache.scala 263:21]
  reg [2:0] value; // @[Counter.scala 29:33]
  wire  _T_87 = io_in_bits_req_cmd == 4'h3; // @[Cache.scala 266:34]
  wire  _T_88 = io_in_bits_req_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_89 = _T_87 | _T_88; // @[Cache.scala 266:62]
  wire  _T_90 = io_out_valid & _T_89; // @[Cache.scala 266:22]
  wire [2:0] _T_93 = value + 3'h1; // @[Counter.scala 39:22]
  wire [2:0] _GEN_0 = _T_90 ? _T_93 : value; // @[Cache.scala 266:85]
  wire  hitWrite = hit & io_in_bits_req_cmd[0]; // @[Cache.scala 270:22]
  wire [63:0] _T_96 = io_in_bits_req_wdata & wordMask; // @[BitUtils.scala 32:13]
  wire [63:0] _T_97 = ~wordMask; // @[BitUtils.scala 32:38]
  wire [63:0] _T_98 = dataRead & _T_97; // @[BitUtils.scala 32:36]
  wire [63:0] dataHitWriteBus_req_bits_data_data = _T_96 | _T_98; // @[BitUtils.scala 32:25]
  wire [2:0] _T_103 = _T_89 ? value : addr_wordIndex; // @[Cache.scala 273:51]
  wire [11:0] dataHitWriteBus_req_bits_setIdx = {addr_index,_T_103}; // @[Cat.scala 29:58]
  wire  _T_105 = ~meta_dirty; // @[Cache.scala 276:25]
  wire  metaHitWriteBus_req_valid = hitWrite & _T_105; // @[Cache.scala 276:22]
  reg [3:0] state; // @[Cache.scala 281:22]
  reg [2:0] value_1; // @[Counter.scala 29:33]
  reg [2:0] value_2; // @[Counter.scala 29:33]
  reg [1:0] state2; // @[Cache.scala 291:23]
  wire  _T_118 = state == 4'h3; // @[Cache.scala 293:39]
  wire  _T_119 = state == 4'h8; // @[Cache.scala 293:66]
  wire  _T_120 = _T_118 | _T_119; // @[Cache.scala 293:57]
  wire  _T_121 = state2 == 2'h0; // @[Cache.scala 293:92]
  wire [2:0] _T_124 = _T_119 ? value_1 : value_2; // @[Cache.scala 294:33]
  wire  _T_126 = state2 == 2'h1; // @[Cache.scala 295:60]
  reg [63:0] dataWay_0_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_1_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_2_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_3_data; // @[Reg.scala 15:16]
  wire [63:0] _T_131 = io_in_bits_waymask[0] ? dataWay_0_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_132 = io_in_bits_waymask[1] ? dataWay_1_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_133 = io_in_bits_waymask[2] ? dataWay_2_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_134 = io_in_bits_waymask[3] ? dataWay_3_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_135 = _T_131 | _T_132; // @[Mux.scala 27:72]
  wire [63:0] _T_136 = _T_135 | _T_133; // @[Mux.scala 27:72]
  wire [63:0] _T_137 = _T_136 | _T_134; // @[Mux.scala 27:72]
  wire  _T_141 = 2'h0 == state2; // @[Conditional.scala 37:30]
  wire  _T_142 = io_dataReadBus_req_ready & io_dataReadBus_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_143 = 2'h1 == state2; // @[Conditional.scala 37:30]
  wire  _T_144 = 2'h2 == state2; // @[Conditional.scala 37:30]
  wire  _T_145 = io_mem_req_ready & io_mem_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_147 = _T_145 | io_cohResp_valid; // @[Cache.scala 301:46]
  wire  _T_149 = _T_147 | hitReadBurst; // @[Cache.scala 301:67]
  wire [31:0] raddr = {io_in_bits_req_addr[31:3],3'h0}; // @[Cat.scala 29:58]
  wire [31:0] waddr = {meta_tag,addr_index,6'h0}; // @[Cat.scala 29:58]
  wire  _T_152 = state == 4'h1; // @[Cache.scala 309:23]
  wire  _T_153 = value_2 == 3'h7; // @[Cache.scala 310:29]
  wire [2:0] _T_154 = _T_153 ? 3'h7 : 3'h3; // @[Cache.scala 310:8]
  wire [2:0] cmd = _T_152 ? 3'h2 : _T_154; // @[Cache.scala 309:16]
  wire  _T_160 = state2 == 2'h2; // @[Cache.scala 316:89]
  wire  _T_161 = _T_118 & _T_160; // @[Cache.scala 316:78]
  reg  afterFirstRead; // @[Cache.scala 323:31]
  reg  alreadyOutFire; // @[Reg.scala 27:20]
  wire  _GEN_12 = io_out_valid | alreadyOutFire; // @[Reg.scala 28:19]
  wire  _T_165 = ~afterFirstRead; // @[Cache.scala 325:22]
  wire  _T_166 = io_mem_resp_ready & io_mem_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_167 = _T_165 & _T_166; // @[Cache.scala 325:38]
  wire  _T_168 = state == 4'h2; // @[Cache.scala 325:70]
  wire  readingFirst = _T_167 & _T_168; // @[Cache.scala 325:60]
  wire  _T_170 = state == 4'h6; // @[Cache.scala 327:52]
  wire  _T_171 = mmio ? _T_170 : readingFirst; // @[Cache.scala 327:39]
  reg [63:0] inRdataRegDemand; // @[Reg.scala 15:16]
  wire  _T_172 = state == 4'h0; // @[Cache.scala 330:31]
  wire  _T_173 = _T_172 & probe; // @[Cache.scala 330:43]
  wire  _T_176 = _T_119 & _T_160; // @[Cache.scala 331:46]
  wire  _T_180 = _T_119 & io_cohResp_valid; // @[Cache.scala 333:49]
  reg [2:0] _T_181; // @[Counter.scala 29:33]
  wire  _T_182 = _T_181 == 3'h7; // @[Counter.scala 38:24]
  wire [2:0] _T_184 = _T_181 + 3'h1; // @[Counter.scala 39:22]
  wire  releaseLast = _T_180 & _T_182; // @[Counter.scala 67:17]
  wire  respToL1Fire = hitReadBurst & _T_160; // @[Cache.scala 337:51]
  wire  _T_195 = _T_172 | _T_176; // @[Cache.scala 338:48]
  wire  _T_196 = _T_195 & hitReadBurst; // @[Cache.scala 338:96]
  reg [2:0] _T_198; // @[Counter.scala 29:33]
  wire  _T_199 = _T_198 == 3'h7; // @[Counter.scala 38:24]
  wire [2:0] _T_201 = _T_198 + 3'h1; // @[Counter.scala 39:22]
  wire  respToL1Last = _T_196 & _T_199; // @[Counter.scala 67:17]
  wire  _T_202 = 4'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_206 = addr_wordIndex == 3'h7; // @[Cache.scala 352:49]
  wire [2:0] _T_208 = addr_wordIndex + 3'h1; // @[Cache.scala 352:93]
  wire  _T_210 = miss | mmio; // @[Cache.scala 353:26]
  wire  _T_217 = 4'h5 == state; // @[Conditional.scala 37:30]
  wire  _T_219 = 4'h6 == state; // @[Conditional.scala 37:30]
  wire  _T_221 = 4'h8 == state; // @[Conditional.scala 37:30]
  wire  _T_223 = io_cohResp_valid | respToL1Fire; // @[Cache.scala 362:31]
  wire [2:0] _T_226 = value_1 + 3'h1; // @[Counter.scala 39:22]
  wire  _T_228 = probe & io_cohResp_valid; // @[Cache.scala 363:19]
  wire  _T_229 = _T_228 & releaseLast; // @[Cache.scala 363:40]
  wire  _T_230 = respToL1Fire & respToL1Last; // @[Cache.scala 363:71]
  wire  _T_231 = _T_229 | _T_230; // @[Cache.scala 363:55]
  wire  _T_232 = 4'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_234 = 4'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_240 = io_mem_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire  _GEN_33 = _T_166 | afterFirstRead; // @[Cache.scala 372:33]
  wire  _T_241 = 4'h3 == state; // @[Conditional.scala 37:30]
  wire [2:0] _T_245 = value_2 + 3'h1; // @[Counter.scala 39:22]
  wire  _T_246 = io_mem_req_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_248 = _T_246 & _T_145; // @[Cache.scala 382:43]
  wire  _T_249 = 4'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_251 = 4'h7 == state; // @[Conditional.scala 37:30]
  wire [63:0] _T_255 = readingFirst ? wordMask : 64'h0; // @[Cache.scala 389:67]
  wire [63:0] _T_256 = io_in_bits_req_wdata & _T_255; // @[BitUtils.scala 32:13]
  wire [63:0] _T_257 = ~_T_255; // @[BitUtils.scala 32:38]
  wire [63:0] _T_258 = io_mem_resp_bits_rdata & _T_257; // @[BitUtils.scala 32:36]
  wire [63:0] dataRefill = _T_256 | _T_258; // @[BitUtils.scala 32:25]
  wire  dataRefillWriteBus_req_valid = _T_168 & _T_166; // @[Cache.scala 391:39]
  wire  metaRefillWriteBus_req_valid = dataRefillWriteBus_req_valid & _T_240; // @[Cache.scala 399:61]
  wire  _T_283 = dataRefillWriteBus_req_valid & _T_8; // @[Cache.scala 409:59]
  wire [2:0] _T_285 = _T_240 ? 3'h6 : 3'h2; // @[Cache.scala 412:29]
  wire  _T_288 = _T_88 | _T_87; // @[Cache.scala 413:35]
  wire [63:0] _T_289 = hit ? dataRead : inRdataRegDemand; // @[Cache.scala 415:31]
  wire  _T_291 = hitReadBurst & _T_119; // @[Cache.scala 417:30]
  wire [2:0] _T_292 = respToL1Last ? 3'h6 : 3'h2; // @[Cache.scala 420:29]
  wire [63:0] _GEN_76 = _T_291 ? _T_137 : _T_289; // @[Cache.scala 417:54]
  wire [3:0] _GEN_77 = _T_291 ? {{1'd0}, _T_292} : io_in_bits_req_cmd; // @[Cache.scala 417:54]
  wire [63:0] _GEN_78 = _T_288 ? _T_289 : _GEN_76; // @[Cache.scala 413:75]
  wire  _T_297 = ~hit; // @[Cache.scala 433:34]
  wire  _T_298 = state == 4'h7; // @[Cache.scala 433:48]
  wire  _T_299 = _T_297 & _T_298; // @[Cache.scala 433:39]
  wire  _T_300 = hit | _T_299; // @[Cache.scala 433:31]
  wire  _T_301 = io_in_bits_req_cmd[0] & _T_300; // @[Cache.scala 433:23]
  wire  _T_307 = _T_301 | _T_283; // @[Cache.scala 433:8]
  wire  _T_310 = _T_230 & _T_119; // @[Cache.scala 433:194]
  wire  _T_311 = _T_307 | _T_310; // @[Cache.scala 433:161]
  wire  _T_313 = io_in_bits_req_cmd[0] | mmio; // @[Cache.scala 434:60]
  wire  _T_315 = ~alreadyOutFire; // @[Cache.scala 434:110]
  wire  _T_316 = afterFirstRead & _T_315; // @[Cache.scala 434:107]
  wire  _T_317 = _T_313 ? _T_298 : _T_316; // @[Cache.scala 434:45]
  wire  _T_318 = hit | _T_317; // @[Cache.scala 434:28]
  wire  _T_319 = probe ? 1'h0 : _T_318; // @[Cache.scala 434:8]
  wire  _T_320 = io_in_bits_req_cmd[1] ? _T_311 : _T_319; // @[Cache.scala 432:37]
  wire  _T_325 = _T_119 & releaseLast; // @[Cache.scala 441:100]
  wire  _T_326 = miss ? _T_172 : _T_325; // @[Cache.scala 441:53]
  wire  _T_327 = io_cohResp_valid & _T_326; // @[Cache.scala 441:47]
  wire  _T_329 = hit | io_in_bits_req_cmd[0]; // @[Cache.scala 442:13]
  wire  _T_334 = _T_298 & _GEN_12; // @[Cache.scala 442:70]
  wire  _T_335 = _T_329 ? io_out_valid : _T_334; // @[Cache.scala 442:8]
  wire  _T_338 = ~hitReadBurst; // @[Cache.scala 445:55]
  wire  _T_339 = _T_172 & _T_338; // @[Cache.scala 445:52]
  wire  _T_341 = ~miss; // @[Cache.scala 445:73]
  wire  _T_342 = _T_339 & _T_341; // @[Cache.scala 445:70]
  wire  _T_343 = ~probe; // @[Cache.scala 445:82]
  wire  _T_352 = metaHitWriteBus_req_valid & metaRefillWriteBus_req_valid; // @[Cache.scala 448:38]
  wire  _T_353 = ~_T_352; // @[Cache.scala 448:10]
  wire  _T_355 = _T_353 | reset; // @[Cache.scala 448:9]
  wire  _T_356 = ~_T_355; // @[Cache.scala 448:9]
  wire  _T_357 = hitWrite & dataRefillWriteBus_req_valid; // @[Cache.scala 449:38]
  wire  _T_358 = ~_T_357; // @[Cache.scala 449:10]
  wire  _T_360 = _T_358 | reset; // @[Cache.scala 449:9]
  wire  _T_361 = ~_T_360; // @[Cache.scala 449:9]
  wire [255:0] _T_376 = {io_in_bits_datas_3_data,io_in_bits_datas_2_data,io_in_bits_datas_1_data,io_in_bits_datas_0_data}; // @[Cache.scala 451:465]
  reg [63:0] _T_377; // @[GTimer.scala 24:20]
  wire [63:0] _T_379 = _T_377 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_383 = ~reset; // @[Debug.scala 56:24]
  reg [63:0] _T_387; // @[GTimer.scala 24:20]
  wire [63:0] _T_389 = _T_387 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_390; // @[GTimer.scala 24:20]
  wire [63:0] _T_392 = _T_390 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_394 = io_metaWriteBus_req_valid & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  reg [63:0] _T_399; // @[GTimer.scala 24:20]
  wire [63:0] _T_401 = _T_399 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_408; // @[GTimer.scala 24:20]
  wire [63:0] _T_410 = _T_408 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_417; // @[GTimer.scala 24:20]
  wire [63:0] _T_419 = _T_417 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_429; // @[GTimer.scala 24:20]
  wire [63:0] _T_431 = _T_429 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_438; // @[GTimer.scala 24:20]
  wire [63:0] _T_440 = _T_438 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_448; // @[GTimer.scala 24:20]
  wire [63:0] _T_450 = _T_448 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_452 = io_dataWriteBus_req_valid & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  wire  _T_459 = _T_118 & _T_145; // @[Cache.scala 460:35]
  reg [63:0] _T_466; // @[GTimer.scala 24:20]
  wire [63:0] _T_468 = _T_466 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_470 = _T_459 & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  wire  _T_477 = _T_152 & _T_145; // @[Cache.scala 461:34]
  reg [63:0] _T_484; // @[GTimer.scala 24:20]
  wire [63:0] _T_486 = _T_484 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_488 = _T_477 & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  reg [63:0] _T_502; // @[GTimer.scala 24:20]
  wire [63:0] _T_504 = _T_502 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_506 = dataRefillWriteBus_req_valid & DISPLAY_ENABLE; // @[Debug.scala 55:16]
  Arbiter_10 metaWriteArb ( // @[Cache.scala 241:28]
    .io_in_0_valid(metaWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(metaWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_tag(metaWriteArb_io_in_0_bits_data_tag),
    .io_in_0_bits_waymask(metaWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(metaWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(metaWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_tag(metaWriteArb_io_in_1_bits_data_tag),
    .io_in_1_bits_data_dirty(metaWriteArb_io_in_1_bits_data_dirty),
    .io_in_1_bits_waymask(metaWriteArb_io_in_1_bits_waymask),
    .io_out_valid(metaWriteArb_io_out_valid),
    .io_out_bits_setIdx(metaWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_tag(metaWriteArb_io_out_bits_data_tag),
    .io_out_bits_data_dirty(metaWriteArb_io_out_bits_data_dirty),
    .io_out_bits_waymask(metaWriteArb_io_out_bits_waymask)
  );
  Arbiter_11 dataWriteArb ( // @[Cache.scala 242:28]
    .io_in_0_valid(dataWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(dataWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_data(dataWriteArb_io_in_0_bits_data_data),
    .io_in_0_bits_waymask(dataWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(dataWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(dataWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_data(dataWriteArb_io_in_1_bits_data_data),
    .io_in_1_bits_waymask(dataWriteArb_io_in_1_bits_waymask),
    .io_out_valid(dataWriteArb_io_out_valid),
    .io_out_bits_setIdx(dataWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_data(dataWriteArb_io_out_bits_data_data),
    .io_out_bits_waymask(dataWriteArb_io_out_bits_waymask)
  );
  assign io_in_ready = _T_342 & _T_343; // @[Cache.scala 445:15]
  assign io_out_valid = io_in_valid & _T_320; // @[Cache.scala 432:16]
  assign io_out_bits_cmd = _T_283 ? {{1'd0}, _T_285} : _GEN_77; // @[Cache.scala 412:23 Cache.scala 420:23 Cache.scala 423:23]
  assign io_out_bits_rdata = _T_283 ? dataRefill : _GEN_78; // @[Cache.scala 411:25 Cache.scala 415:25 Cache.scala 419:25 Cache.scala 422:25]
  assign io_isFinish = probe ? _T_327 : _T_335; // @[Cache.scala 441:15]
  assign io_dataReadBus_req_valid = _T_120 & _T_121; // @[SRAMTemplate.scala 53:20]
  assign io_dataReadBus_req_bits_setIdx = {addr_index,_T_124}; // @[SRAMTemplate.scala 26:17]
  assign io_dataWriteBus_req_valid = dataWriteArb_io_out_valid; // @[Cache.scala 396:23]
  assign io_dataWriteBus_req_bits_setIdx = dataWriteArb_io_out_bits_setIdx; // @[Cache.scala 396:23]
  assign io_dataWriteBus_req_bits_data_data = dataWriteArb_io_out_bits_data_data; // @[Cache.scala 396:23]
  assign io_dataWriteBus_req_bits_waymask = dataWriteArb_io_out_bits_waymask; // @[Cache.scala 396:23]
  assign io_metaWriteBus_req_valid = metaWriteArb_io_out_valid; // @[Cache.scala 406:23]
  assign io_metaWriteBus_req_bits_setIdx = metaWriteArb_io_out_bits_setIdx; // @[Cache.scala 406:23]
  assign io_metaWriteBus_req_bits_data_tag = metaWriteArb_io_out_bits_data_tag; // @[Cache.scala 406:23]
  assign io_metaWriteBus_req_bits_data_valid = 1'h1; // @[Cache.scala 406:23]
  assign io_metaWriteBus_req_bits_data_dirty = metaWriteArb_io_out_bits_data_dirty; // @[Cache.scala 406:23]
  assign io_metaWriteBus_req_bits_waymask = metaWriteArb_io_out_bits_waymask; // @[Cache.scala 406:23]
  assign io_mem_req_valid = _T_152 | _T_161; // @[Cache.scala 316:20]
  assign io_mem_req_bits_addr = _T_152 ? raddr : waddr; // @[SimpleBus.scala 64:15]
  assign io_mem_req_bits_size = 3'h3; // @[SimpleBus.scala 66:15]
  assign io_mem_req_bits_cmd = {{1'd0}, cmd}; // @[SimpleBus.scala 65:14]
  assign io_mem_req_bits_wmask = 8'hff; // @[SimpleBus.scala 68:16]
  assign io_mem_req_bits_wdata = _T_136 | _T_134; // @[SimpleBus.scala 67:16]
  assign io_mem_resp_ready = 1'h1; // @[Cache.scala 315:21]
  assign io_cohResp_valid = _T_173 | _T_176; // @[Cache.scala 330:20]
  assign io_dataReadRespToL1 = hitReadBurst & _T_195; // @[Cache.scala 446:23]
  assign metaWriteArb_io_in_0_valid = hitWrite & _T_105; // @[Cache.scala 404:25]
  assign metaWriteArb_io_in_0_bits_setIdx = io_in_bits_req_addr[14:6]; // @[Cache.scala 404:25]
  assign metaWriteArb_io_in_0_bits_data_tag = _T_27[18:2]; // @[Cache.scala 404:25]
  assign metaWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[Cache.scala 404:25]
  assign metaWriteArb_io_in_1_valid = dataRefillWriteBus_req_valid & _T_240; // @[Cache.scala 405:25]
  assign metaWriteArb_io_in_1_bits_setIdx = io_in_bits_req_addr[14:6]; // @[Cache.scala 405:25]
  assign metaWriteArb_io_in_1_bits_data_tag = io_in_bits_req_addr[31:15]; // @[Cache.scala 405:25]
  assign metaWriteArb_io_in_1_bits_data_dirty = io_in_bits_req_cmd[0]; // @[Cache.scala 405:25]
  assign metaWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[Cache.scala 405:25]
  assign dataWriteArb_io_in_0_valid = hit & io_in_bits_req_cmd[0]; // @[Cache.scala 394:25]
  assign dataWriteArb_io_in_0_bits_setIdx = {addr_index,_T_103}; // @[Cache.scala 394:25]
  assign dataWriteArb_io_in_0_bits_data_data = _T_96 | _T_98; // @[Cache.scala 394:25]
  assign dataWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[Cache.scala 394:25]
  assign dataWriteArb_io_in_1_valid = _T_168 & _T_166; // @[Cache.scala 395:25]
  assign dataWriteArb_io_in_1_bits_setIdx = {addr_index,value_1}; // @[Cache.scala 395:25]
  assign dataWriteArb_io_in_1_bits_data_data = _T_256 | _T_258; // @[Cache.scala 395:25]
  assign dataWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[Cache.scala 395:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  value_2 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  state2 = _RAND_4[1:0];
  _RAND_5 = {2{`RANDOM}};
  dataWay_0_data = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  dataWay_1_data = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  dataWay_2_data = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  dataWay_3_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  afterFirstRead = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  alreadyOutFire = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  inRdataRegDemand = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  _T_181 = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  _T_198 = _RAND_13[2:0];
  _RAND_14 = {2{`RANDOM}};
  _T_377 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  _T_387 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  _T_390 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  _T_399 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  _T_408 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  _T_417 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  _T_429 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  _T_438 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  _T_448 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  _T_466 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  _T_484 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  _T_502 = _RAND_25[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 3'h0;
    end else if (_T_202) begin
      if (_T_90) begin
        value <= _T_93;
      end
    end else if (_T_217) begin
      if (_T_90) begin
        value <= _T_93;
      end
    end else if (_T_219) begin
      if (_T_90) begin
        value <= _T_93;
      end
    end else if (_T_221) begin
      if (_T_90) begin
        value <= _T_93;
      end
    end else if (_T_232) begin
      value <= _GEN_0;
    end else if (_T_234) begin
      if (_T_166) begin
        if (_T_87) begin
          value <= 3'h0;
        end else begin
          value <= _GEN_0;
        end
      end else begin
        value <= _GEN_0;
      end
    end else begin
      value <= _GEN_0;
    end
    if (reset) begin
      state <= 4'h0;
    end else if (_T_202) begin
      if (probe) begin
        if (io_cohResp_valid) begin
          if (hit) begin
            state <= 4'h8;
          end else begin
            state <= 4'h0;
          end
        end
      end else if (hitReadBurst) begin
        state <= 4'h8;
      end else if (_T_210) begin
        if (mmio) begin
          state <= 4'h5;
        end else if (meta_dirty) begin
          state <= 4'h3;
        end else begin
          state <= 4'h1;
        end
      end
    end else if (!(_T_217)) begin
      if (!(_T_219)) begin
        if (_T_221) begin
          if (_T_231) begin
            state <= 4'h0;
          end
        end else if (_T_232) begin
          if (_T_145) begin
            state <= 4'h2;
          end
        end else if (_T_234) begin
          if (_T_166) begin
            if (_T_240) begin
              state <= 4'h7;
            end
          end
        end else if (_T_241) begin
          if (_T_248) begin
            state <= 4'h4;
          end
        end else if (_T_249) begin
          if (_T_166) begin
            state <= 4'h1;
          end
        end else if (_T_251) begin
          if (_GEN_12) begin
            state <= 4'h0;
          end
        end
      end
    end
    if (reset) begin
      value_1 <= 3'h0;
    end else if (_T_202) begin
      if (probe) begin
        if (io_cohResp_valid) begin
          value_1 <= addr_wordIndex;
        end
      end else if (hitReadBurst) begin
        if (_T_206) begin
          value_1 <= 3'h0;
        end else begin
          value_1 <= _T_208;
        end
      end
    end else if (!(_T_217)) begin
      if (!(_T_219)) begin
        if (_T_221) begin
          if (_T_223) begin
            value_1 <= _T_226;
          end
        end else if (_T_232) begin
          if (_T_145) begin
            value_1 <= addr_wordIndex;
          end
        end else if (_T_234) begin
          if (_T_166) begin
            value_1 <= _T_226;
          end
        end
      end
    end
    if (reset) begin
      value_2 <= 3'h0;
    end else if (!(_T_202)) begin
      if (!(_T_217)) begin
        if (!(_T_219)) begin
          if (!(_T_221)) begin
            if (!(_T_232)) begin
              if (!(_T_234)) begin
                if (_T_241) begin
                  if (_T_145) begin
                    value_2 <= _T_245;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      state2 <= 2'h0;
    end else if (_T_141) begin
      if (_T_142) begin
        state2 <= 2'h1;
      end
    end else if (_T_143) begin
      state2 <= 2'h2;
    end else if (_T_144) begin
      if (_T_149) begin
        state2 <= 2'h0;
      end
    end
    if (_T_126) begin
      dataWay_0_data <= io_dataReadBus_resp_data_0_data;
    end
    if (_T_126) begin
      dataWay_1_data <= io_dataReadBus_resp_data_1_data;
    end
    if (_T_126) begin
      dataWay_2_data <= io_dataReadBus_resp_data_2_data;
    end
    if (_T_126) begin
      dataWay_3_data <= io_dataReadBus_resp_data_3_data;
    end
    if (reset) begin
      afterFirstRead <= 1'h0;
    end else if (_T_202) begin
      afterFirstRead <= 1'h0;
    end else if (!(_T_217)) begin
      if (!(_T_219)) begin
        if (!(_T_221)) begin
          if (!(_T_232)) begin
            if (_T_234) begin
              afterFirstRead <= _GEN_33;
            end
          end
        end
      end
    end
    if (reset) begin
      alreadyOutFire <= 1'h0;
    end else if (_T_202) begin
      alreadyOutFire <= 1'h0;
    end else begin
      alreadyOutFire <= _GEN_12;
    end
    if (_T_171) begin
      if (mmio) begin
        inRdataRegDemand <= 64'h0;
      end else begin
        inRdataRegDemand <= io_mem_resp_bits_rdata;
      end
    end
    if (reset) begin
      _T_181 <= 3'h0;
    end else if (_T_180) begin
      _T_181 <= _T_184;
    end
    if (reset) begin
      _T_198 <= 3'h0;
    end else if (_T_196) begin
      _T_198 <= _T_201;
    end
    if (reset) begin
      _T_377 <= 64'h0;
    end else begin
      _T_377 <= _T_379;
    end
    if (reset) begin
      _T_387 <= 64'h0;
    end else begin
      _T_387 <= _T_389;
    end
    if (reset) begin
      _T_390 <= 64'h0;
    end else begin
      _T_390 <= _T_392;
    end
    if (reset) begin
      _T_399 <= 64'h0;
    end else begin
      _T_399 <= _T_401;
    end
    if (reset) begin
      _T_408 <= 64'h0;
    end else begin
      _T_408 <= _T_410;
    end
    if (reset) begin
      _T_417 <= 64'h0;
    end else begin
      _T_417 <= _T_419;
    end
    if (reset) begin
      _T_429 <= 64'h0;
    end else begin
      _T_429 <= _T_431;
    end
    if (reset) begin
      _T_438 <= 64'h0;
    end else begin
      _T_438 <= _T_440;
    end
    if (reset) begin
      _T_448 <= 64'h0;
    end else begin
      _T_448 <= _T_450;
    end
    if (reset) begin
      _T_466 <= 64'h0;
    end else begin
      _T_466 <= _T_468;
    end
    if (reset) begin
      _T_484 <= 64'h0;
    end else begin
      _T_484 <= _T_486;
    end
    if (reset) begin
      _T_502 <= 64'h0;
    end else begin
      _T_502 <= _T_504;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_36) begin
          $fwrite(32'h80000002,"Assertion failed: MMIO request should not hit in cache\n    at Cache.scala:252 assert(!(mmio && hit), \"MMIO request should not hit in cache\")\n"); // @[Cache.scala 252:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_36) begin
          $fatal; // @[Cache.scala 252:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_356) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Cache.scala:448 assert(!(metaHitWriteBus.req.valid && metaRefillWriteBus.req.valid))\n"); // @[Cache.scala 448:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_356) begin
          $fatal; // @[Cache.scala 448:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_361) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Cache.scala:449 assert(!(dataHitWriteBus.req.valid && dataRefillWriteBus.req.valid))\n"); // @[Cache.scala 449:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_361) begin
          $fatal; // @[Cache.scala 449:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_383) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_2: ",_T_377); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_383) begin
          $fwrite(32'h80000002," metaread idx %x waymask %b metas %x%x:%x %x%x:%x %x%x:%x %x%x:%x %x\n",addr_index,io_in_bits_waymask,io_in_bits_metas_0_valid,io_in_bits_metas_0_dirty,io_in_bits_metas_0_tag,io_in_bits_metas_1_valid,io_in_bits_metas_1_dirty,io_in_bits_metas_1_tag,io_in_bits_metas_2_valid,io_in_bits_metas_2_dirty,io_in_bits_metas_2_tag,io_in_bits_metas_3_valid,io_in_bits_metas_3_dirty,io_in_bits_metas_3_tag,_T_376); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_394 & _T_383) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_2: ",_T_390); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_394 & _T_383) begin
          $fwrite(32'h80000002,"%d: [l2cache S3]: metawrite idx %x wmask %b meta %x%x:%x\n",_T_387,io_metaWriteBus_req_bits_setIdx,io_metaWriteBus_req_bits_waymask,io_metaWriteBus_req_bits_data_valid,io_metaWriteBus_req_bits_data_dirty,io_metaWriteBus_req_bits_data_tag); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_383) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_2: ",_T_399); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_383) begin
          $fwrite(32'h80000002," in.ready = %d, in.valid = %d, hit = %x, state = %d, addr = %x cmd:%d probe:%d isFinish:%d\n",io_in_ready,io_in_valid,hit,state,io_in_bits_req_addr,io_in_bits_req_cmd,probe,io_isFinish); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_383) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_2: ",_T_408); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_383) begin
          $fwrite(32'h80000002," out.valid:%d rdata:%x cmd:%d user:%x id:%x \n",io_out_valid,io_out_bits_rdata,io_out_bits_cmd,1'h0,1'h0); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_383) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_2: ",_T_417); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_383) begin
          $fwrite(32'h80000002," DHW: (%d, %d), data:%x setIdx:%x MHW:(%d, %d)\n",hitWrite,1'h1,dataHitWriteBus_req_bits_data_data,dataHitWriteBus_req_bits_setIdx,metaHitWriteBus_req_valid,1'h1); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_383) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_2: ",_T_429); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_383) begin
          $fwrite(32'h80000002," DreadCache: %x \n",_T_376); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_383) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_2: ",_T_438); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_383) begin
          $fwrite(32'h80000002," useFD:%d isFD:%d FD:%x DreadArray:%x dataRead:%x inwaymask:%x FDwaymask:%x \n",useForwardData,io_in_bits_isForwardData,io_in_bits_forwardData_data_data,_T_48,dataRead,io_in_bits_waymask,io_in_bits_forwardData_waymask); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_452 & _T_383) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_2: ",_T_448); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_452 & _T_383) begin
          $fwrite(32'h80000002,"[WB] waymask: %b data:%x setIdx:%x\n",io_dataWriteBus_req_bits_waymask,io_dataWriteBus_req_bits_data_data,io_dataWriteBus_req_bits_setIdx); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_470 & _T_383) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_2: ",_T_466); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_470 & _T_383) begin
          $fwrite(32'h80000002,"[COUTW] cnt %x addr %x data %x cmd %x size %x wmask %x tag %x idx %x waymask %b \n",value_2,io_mem_req_bits_addr,io_mem_req_bits_wdata,io_mem_req_bits_cmd,io_mem_req_bits_size,io_mem_req_bits_wmask,addr_tag,addr_index,io_in_bits_waymask); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_488 & _T_383) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_2: ",_T_484); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_488 & _T_383) begin
          $fwrite(32'h80000002,"[COUTR] addr %x tag %x idx %x waymask %b \n",io_mem_req_bits_addr,addr_tag,addr_index,io_in_bits_waymask); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_506 & _T_383) begin
          $fwrite(32'h80000002,"[%d] CacheStage3_2: ",_T_502); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_506 & _T_383) begin
          $fwrite(32'h80000002,"[COUTR] cnt %x data %x tag %x idx %x waymask %b \n",value_1,io_mem_resp_bits_rdata,addr_tag,addr_index,io_in_bits_waymask); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module SRAMTemplate_5(
  input         clock,
  input         reset,
  output        io_r_req_ready,
  input         io_r_req_valid,
  input  [8:0]  io_r_req_bits_setIdx,
  output [16:0] io_r_resp_data_0_tag,
  output        io_r_resp_data_0_valid,
  output        io_r_resp_data_0_dirty,
  output [16:0] io_r_resp_data_1_tag,
  output        io_r_resp_data_1_valid,
  output        io_r_resp_data_1_dirty,
  output [16:0] io_r_resp_data_2_tag,
  output        io_r_resp_data_2_valid,
  output        io_r_resp_data_2_dirty,
  output [16:0] io_r_resp_data_3_tag,
  output        io_r_resp_data_3_valid,
  output        io_r_resp_data_3_dirty,
  input         io_w_req_valid,
  input  [8:0]  io_w_req_bits_setIdx,
  input  [16:0] io_w_req_bits_data_tag,
  input         io_w_req_bits_data_dirty,
  input  [3:0]  io_w_req_bits_waymask
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  reg [18:0] array_0 [0:511]; // @[SRAMTemplate.scala 76:26]
  wire [18:0] array_0__T_21_data; // @[SRAMTemplate.scala 76:26]
  wire [8:0] array_0__T_21_addr; // @[SRAMTemplate.scala 76:26]
  wire [18:0] array_0__T_17_data; // @[SRAMTemplate.scala 76:26]
  wire [8:0] array_0__T_17_addr; // @[SRAMTemplate.scala 76:26]
  wire  array_0__T_17_mask; // @[SRAMTemplate.scala 76:26]
  wire  array_0__T_17_en; // @[SRAMTemplate.scala 76:26]
  reg  array_0__T_21_en_pipe_0;
  reg [8:0] array_0__T_21_addr_pipe_0;
  reg [18:0] array_1 [0:511]; // @[SRAMTemplate.scala 76:26]
  wire [18:0] array_1__T_21_data; // @[SRAMTemplate.scala 76:26]
  wire [8:0] array_1__T_21_addr; // @[SRAMTemplate.scala 76:26]
  wire [18:0] array_1__T_17_data; // @[SRAMTemplate.scala 76:26]
  wire [8:0] array_1__T_17_addr; // @[SRAMTemplate.scala 76:26]
  wire  array_1__T_17_mask; // @[SRAMTemplate.scala 76:26]
  wire  array_1__T_17_en; // @[SRAMTemplate.scala 76:26]
  reg  array_1__T_21_en_pipe_0;
  reg [8:0] array_1__T_21_addr_pipe_0;
  reg [18:0] array_2 [0:511]; // @[SRAMTemplate.scala 76:26]
  wire [18:0] array_2__T_21_data; // @[SRAMTemplate.scala 76:26]
  wire [8:0] array_2__T_21_addr; // @[SRAMTemplate.scala 76:26]
  wire [18:0] array_2__T_17_data; // @[SRAMTemplate.scala 76:26]
  wire [8:0] array_2__T_17_addr; // @[SRAMTemplate.scala 76:26]
  wire  array_2__T_17_mask; // @[SRAMTemplate.scala 76:26]
  wire  array_2__T_17_en; // @[SRAMTemplate.scala 76:26]
  reg  array_2__T_21_en_pipe_0;
  reg [8:0] array_2__T_21_addr_pipe_0;
  reg [18:0] array_3 [0:511]; // @[SRAMTemplate.scala 76:26]
  wire [18:0] array_3__T_21_data; // @[SRAMTemplate.scala 76:26]
  wire [8:0] array_3__T_21_addr; // @[SRAMTemplate.scala 76:26]
  wire [18:0] array_3__T_17_data; // @[SRAMTemplate.scala 76:26]
  wire [8:0] array_3__T_17_addr; // @[SRAMTemplate.scala 76:26]
  wire  array_3__T_17_mask; // @[SRAMTemplate.scala 76:26]
  wire  array_3__T_17_en; // @[SRAMTemplate.scala 76:26]
  reg  array_3__T_21_en_pipe_0;
  reg [8:0] array_3__T_21_addr_pipe_0;
  reg  resetState; // @[SRAMTemplate.scala 80:30]
  reg [8:0] resetSet; // @[Counter.scala 29:33]
  wire  _T_3 = resetSet == 9'h1ff; // @[Counter.scala 38:24]
  wire [8:0] _T_5 = resetSet + 9'h1; // @[Counter.scala 39:22]
  wire  _GEN_1 = resetState & _T_3; // @[Counter.scala 67:17]
  wire  _GEN_2 = _GEN_1 ? 1'h0 : resetState; // @[SRAMTemplate.scala 82:24]
  wire  wen = io_w_req_valid | resetState; // @[SRAMTemplate.scala 88:52]
  wire  _T_6 = ~wen; // @[SRAMTemplate.scala 89:41]
  wire [18:0] _T_9 = {io_w_req_bits_data_tag,1'h1,io_w_req_bits_data_dirty}; // @[SRAMTemplate.scala 92:78]
  wire [3:0] waymask = resetState ? 4'hf : io_w_req_bits_waymask; // @[SRAMTemplate.scala 93:20]
  wire [18:0] _T_22 = array_0__T_21_data;
  wire [18:0] _T_26 = array_1__T_21_data;
  wire [18:0] _T_30 = array_2__T_21_data;
  wire [18:0] _T_34 = array_3__T_21_data;
  wire  _T_39 = ~resetState; // @[SRAMTemplate.scala 101:21]
  assign array_0__T_21_addr = array_0__T_21_addr_pipe_0;
  assign array_0__T_21_data = array_0[array_0__T_21_addr]; // @[SRAMTemplate.scala 76:26]
  assign array_0__T_17_data = resetState ? 19'h0 : _T_9;
  assign array_0__T_17_addr = resetState ? resetSet : io_w_req_bits_setIdx;
  assign array_0__T_17_mask = waymask[0];
  assign array_0__T_17_en = io_w_req_valid | resetState;
  assign array_1__T_21_addr = array_1__T_21_addr_pipe_0;
  assign array_1__T_21_data = array_1[array_1__T_21_addr]; // @[SRAMTemplate.scala 76:26]
  assign array_1__T_17_data = resetState ? 19'h0 : _T_9;
  assign array_1__T_17_addr = resetState ? resetSet : io_w_req_bits_setIdx;
  assign array_1__T_17_mask = waymask[1];
  assign array_1__T_17_en = io_w_req_valid | resetState;
  assign array_2__T_21_addr = array_2__T_21_addr_pipe_0;
  assign array_2__T_21_data = array_2[array_2__T_21_addr]; // @[SRAMTemplate.scala 76:26]
  assign array_2__T_17_data = resetState ? 19'h0 : _T_9;
  assign array_2__T_17_addr = resetState ? resetSet : io_w_req_bits_setIdx;
  assign array_2__T_17_mask = waymask[2];
  assign array_2__T_17_en = io_w_req_valid | resetState;
  assign array_3__T_21_addr = array_3__T_21_addr_pipe_0;
  assign array_3__T_21_data = array_3[array_3__T_21_addr]; // @[SRAMTemplate.scala 76:26]
  assign array_3__T_17_data = resetState ? 19'h0 : _T_9;
  assign array_3__T_17_addr = resetState ? resetSet : io_w_req_bits_setIdx;
  assign array_3__T_17_mask = waymask[3];
  assign array_3__T_17_en = io_w_req_valid | resetState;
  assign io_r_req_ready = _T_39 & _T_6; // @[SRAMTemplate.scala 101:18]
  assign io_r_resp_data_0_tag = _T_22[18:2]; // @[SRAMTemplate.scala 99:18]
  assign io_r_resp_data_0_valid = _T_22[1]; // @[SRAMTemplate.scala 99:18]
  assign io_r_resp_data_0_dirty = _T_22[0]; // @[SRAMTemplate.scala 99:18]
  assign io_r_resp_data_1_tag = _T_26[18:2]; // @[SRAMTemplate.scala 99:18]
  assign io_r_resp_data_1_valid = _T_26[1]; // @[SRAMTemplate.scala 99:18]
  assign io_r_resp_data_1_dirty = _T_26[0]; // @[SRAMTemplate.scala 99:18]
  assign io_r_resp_data_2_tag = _T_30[18:2]; // @[SRAMTemplate.scala 99:18]
  assign io_r_resp_data_2_valid = _T_30[1]; // @[SRAMTemplate.scala 99:18]
  assign io_r_resp_data_2_dirty = _T_30[0]; // @[SRAMTemplate.scala 99:18]
  assign io_r_resp_data_3_tag = _T_34[18:2]; // @[SRAMTemplate.scala 99:18]
  assign io_r_resp_data_3_valid = _T_34[1]; // @[SRAMTemplate.scala 99:18]
  assign io_r_resp_data_3_dirty = _T_34[0]; // @[SRAMTemplate.scala 99:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    array_0[initvar] = _RAND_0[18:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    array_1[initvar] = _RAND_3[18:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    array_2[initvar] = _RAND_6[18:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    array_3[initvar] = _RAND_9[18:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  array_0__T_21_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  array_0__T_21_addr_pipe_0 = _RAND_2[8:0];
  _RAND_4 = {1{`RANDOM}};
  array_1__T_21_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  array_1__T_21_addr_pipe_0 = _RAND_5[8:0];
  _RAND_7 = {1{`RANDOM}};
  array_2__T_21_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  array_2__T_21_addr_pipe_0 = _RAND_8[8:0];
  _RAND_10 = {1{`RANDOM}};
  array_3__T_21_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  array_3__T_21_addr_pipe_0 = _RAND_11[8:0];
  _RAND_12 = {1{`RANDOM}};
  resetState = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  resetSet = _RAND_13[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(array_0__T_17_en & array_0__T_17_mask) begin
      array_0[array_0__T_17_addr] <= array_0__T_17_data; // @[SRAMTemplate.scala 76:26]
    end
    array_0__T_21_en_pipe_0 <= io_r_req_valid & _T_6;
    if (io_r_req_valid & _T_6) begin
      array_0__T_21_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if(array_1__T_17_en & array_1__T_17_mask) begin
      array_1[array_1__T_17_addr] <= array_1__T_17_data; // @[SRAMTemplate.scala 76:26]
    end
    array_1__T_21_en_pipe_0 <= io_r_req_valid & _T_6;
    if (io_r_req_valid & _T_6) begin
      array_1__T_21_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if(array_2__T_17_en & array_2__T_17_mask) begin
      array_2[array_2__T_17_addr] <= array_2__T_17_data; // @[SRAMTemplate.scala 76:26]
    end
    array_2__T_21_en_pipe_0 <= io_r_req_valid & _T_6;
    if (io_r_req_valid & _T_6) begin
      array_2__T_21_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if(array_3__T_17_en & array_3__T_17_mask) begin
      array_3[array_3__T_17_addr] <= array_3__T_17_data; // @[SRAMTemplate.scala 76:26]
    end
    array_3__T_21_en_pipe_0 <= io_r_req_valid & _T_6;
    if (io_r_req_valid & _T_6) begin
      array_3__T_21_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    resetState <= reset | _GEN_2;
    if (reset) begin
      resetSet <= 9'h0;
    end else if (resetState) begin
      resetSet <= _T_5;
    end
  end
endmodule
module Arbiter_12(
  output       io_in_0_ready,
  input        io_in_0_valid,
  input  [8:0] io_in_0_bits_setIdx,
  input        io_out_ready,
  output       io_out_valid,
  output [8:0] io_out_bits_setIdx
);
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:14]
  assign io_out_valid = io_in_0_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_setIdx = io_in_0_bits_setIdx; // @[Arbiter.scala 124:15]
endmodule
module SRAMTemplateWithArbiter_4(
  input         clock,
  input         reset,
  output        io_r_0_req_ready,
  input         io_r_0_req_valid,
  input  [8:0]  io_r_0_req_bits_setIdx,
  output [16:0] io_r_0_resp_data_0_tag,
  output        io_r_0_resp_data_0_valid,
  output        io_r_0_resp_data_0_dirty,
  output [16:0] io_r_0_resp_data_1_tag,
  output        io_r_0_resp_data_1_valid,
  output        io_r_0_resp_data_1_dirty,
  output [16:0] io_r_0_resp_data_2_tag,
  output        io_r_0_resp_data_2_valid,
  output        io_r_0_resp_data_2_dirty,
  output [16:0] io_r_0_resp_data_3_tag,
  output        io_r_0_resp_data_3_valid,
  output        io_r_0_resp_data_3_dirty,
  input         io_w_req_valid,
  input  [8:0]  io_w_req_bits_setIdx,
  input  [16:0] io_w_req_bits_data_tag,
  input         io_w_req_bits_data_dirty,
  input  [3:0]  io_w_req_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  ram_clock; // @[SRAMTemplate.scala 121:19]
  wire  ram_reset; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_r_req_ready; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_r_req_valid; // @[SRAMTemplate.scala 121:19]
  wire [8:0] ram_io_r_req_bits_setIdx; // @[SRAMTemplate.scala 121:19]
  wire [16:0] ram_io_r_resp_data_0_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_r_resp_data_0_valid; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_r_resp_data_0_dirty; // @[SRAMTemplate.scala 121:19]
  wire [16:0] ram_io_r_resp_data_1_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_r_resp_data_1_valid; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_r_resp_data_1_dirty; // @[SRAMTemplate.scala 121:19]
  wire [16:0] ram_io_r_resp_data_2_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_r_resp_data_2_valid; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_r_resp_data_2_dirty; // @[SRAMTemplate.scala 121:19]
  wire [16:0] ram_io_r_resp_data_3_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_r_resp_data_3_valid; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_r_resp_data_3_dirty; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_w_req_valid; // @[SRAMTemplate.scala 121:19]
  wire [8:0] ram_io_w_req_bits_setIdx; // @[SRAMTemplate.scala 121:19]
  wire [16:0] ram_io_w_req_bits_data_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_w_req_bits_data_dirty; // @[SRAMTemplate.scala 121:19]
  wire [3:0] ram_io_w_req_bits_waymask; // @[SRAMTemplate.scala 121:19]
  wire  readArb_io_in_0_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_in_0_valid; // @[SRAMTemplate.scala 124:23]
  wire [8:0] readArb_io_in_0_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_out_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_out_valid; // @[SRAMTemplate.scala 124:23]
  wire [8:0] readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  reg  _T_1; // @[SRAMTemplate.scala 130:58]
  reg [16:0] _T_3_0_tag; // @[Reg.scala 27:20]
  reg  _T_3_0_valid; // @[Reg.scala 27:20]
  reg  _T_3_0_dirty; // @[Reg.scala 27:20]
  reg [16:0] _T_3_1_tag; // @[Reg.scala 27:20]
  reg  _T_3_1_valid; // @[Reg.scala 27:20]
  reg  _T_3_1_dirty; // @[Reg.scala 27:20]
  reg [16:0] _T_3_2_tag; // @[Reg.scala 27:20]
  reg  _T_3_2_valid; // @[Reg.scala 27:20]
  reg  _T_3_2_dirty; // @[Reg.scala 27:20]
  reg [16:0] _T_3_3_tag; // @[Reg.scala 27:20]
  reg  _T_3_3_valid; // @[Reg.scala 27:20]
  reg  _T_3_3_dirty; // @[Reg.scala 27:20]
  SRAMTemplate_5 ram ( // @[SRAMTemplate.scala 121:19]
    .clock(ram_clock),
    .reset(ram_reset),
    .io_r_req_ready(ram_io_r_req_ready),
    .io_r_req_valid(ram_io_r_req_valid),
    .io_r_req_bits_setIdx(ram_io_r_req_bits_setIdx),
    .io_r_resp_data_0_tag(ram_io_r_resp_data_0_tag),
    .io_r_resp_data_0_valid(ram_io_r_resp_data_0_valid),
    .io_r_resp_data_0_dirty(ram_io_r_resp_data_0_dirty),
    .io_r_resp_data_1_tag(ram_io_r_resp_data_1_tag),
    .io_r_resp_data_1_valid(ram_io_r_resp_data_1_valid),
    .io_r_resp_data_1_dirty(ram_io_r_resp_data_1_dirty),
    .io_r_resp_data_2_tag(ram_io_r_resp_data_2_tag),
    .io_r_resp_data_2_valid(ram_io_r_resp_data_2_valid),
    .io_r_resp_data_2_dirty(ram_io_r_resp_data_2_dirty),
    .io_r_resp_data_3_tag(ram_io_r_resp_data_3_tag),
    .io_r_resp_data_3_valid(ram_io_r_resp_data_3_valid),
    .io_r_resp_data_3_dirty(ram_io_r_resp_data_3_dirty),
    .io_w_req_valid(ram_io_w_req_valid),
    .io_w_req_bits_setIdx(ram_io_w_req_bits_setIdx),
    .io_w_req_bits_data_tag(ram_io_w_req_bits_data_tag),
    .io_w_req_bits_data_dirty(ram_io_w_req_bits_data_dirty),
    .io_w_req_bits_waymask(ram_io_w_req_bits_waymask)
  );
  Arbiter_12 readArb ( // @[SRAMTemplate.scala 124:23]
    .io_in_0_ready(readArb_io_in_0_ready),
    .io_in_0_valid(readArb_io_in_0_valid),
    .io_in_0_bits_setIdx(readArb_io_in_0_bits_setIdx),
    .io_out_ready(readArb_io_out_ready),
    .io_out_valid(readArb_io_out_valid),
    .io_out_bits_setIdx(readArb_io_out_bits_setIdx)
  );
  assign io_r_0_req_ready = readArb_io_in_0_ready; // @[SRAMTemplate.scala 125:17]
  assign io_r_0_resp_data_0_tag = _T_1 ? ram_io_r_resp_data_0_tag : _T_3_0_tag; // @[SRAMTemplate.scala 130:17]
  assign io_r_0_resp_data_0_valid = _T_1 ? ram_io_r_resp_data_0_valid : _T_3_0_valid; // @[SRAMTemplate.scala 130:17]
  assign io_r_0_resp_data_0_dirty = _T_1 ? ram_io_r_resp_data_0_dirty : _T_3_0_dirty; // @[SRAMTemplate.scala 130:17]
  assign io_r_0_resp_data_1_tag = _T_1 ? ram_io_r_resp_data_1_tag : _T_3_1_tag; // @[SRAMTemplate.scala 130:17]
  assign io_r_0_resp_data_1_valid = _T_1 ? ram_io_r_resp_data_1_valid : _T_3_1_valid; // @[SRAMTemplate.scala 130:17]
  assign io_r_0_resp_data_1_dirty = _T_1 ? ram_io_r_resp_data_1_dirty : _T_3_1_dirty; // @[SRAMTemplate.scala 130:17]
  assign io_r_0_resp_data_2_tag = _T_1 ? ram_io_r_resp_data_2_tag : _T_3_2_tag; // @[SRAMTemplate.scala 130:17]
  assign io_r_0_resp_data_2_valid = _T_1 ? ram_io_r_resp_data_2_valid : _T_3_2_valid; // @[SRAMTemplate.scala 130:17]
  assign io_r_0_resp_data_2_dirty = _T_1 ? ram_io_r_resp_data_2_dirty : _T_3_2_dirty; // @[SRAMTemplate.scala 130:17]
  assign io_r_0_resp_data_3_tag = _T_1 ? ram_io_r_resp_data_3_tag : _T_3_3_tag; // @[SRAMTemplate.scala 130:17]
  assign io_r_0_resp_data_3_valid = _T_1 ? ram_io_r_resp_data_3_valid : _T_3_3_valid; // @[SRAMTemplate.scala 130:17]
  assign io_r_0_resp_data_3_dirty = _T_1 ? ram_io_r_resp_data_3_dirty : _T_3_3_dirty; // @[SRAMTemplate.scala 130:17]
  assign ram_clock = clock;
  assign ram_reset = reset;
  assign ram_io_r_req_valid = readArb_io_out_valid; // @[SRAMTemplate.scala 126:16]
  assign ram_io_r_req_bits_setIdx = readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 126:16]
  assign ram_io_w_req_valid = io_w_req_valid; // @[SRAMTemplate.scala 122:12]
  assign ram_io_w_req_bits_setIdx = io_w_req_bits_setIdx; // @[SRAMTemplate.scala 122:12]
  assign ram_io_w_req_bits_data_tag = io_w_req_bits_data_tag; // @[SRAMTemplate.scala 122:12]
  assign ram_io_w_req_bits_data_dirty = io_w_req_bits_data_dirty; // @[SRAMTemplate.scala 122:12]
  assign ram_io_w_req_bits_waymask = io_w_req_bits_waymask; // @[SRAMTemplate.scala 122:12]
  assign readArb_io_in_0_valid = io_r_0_req_valid; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_in_0_bits_setIdx = io_r_0_req_bits_setIdx; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_out_ready = ram_io_r_req_ready; // @[SRAMTemplate.scala 126:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _T_3_0_tag = _RAND_1[16:0];
  _RAND_2 = {1{`RANDOM}};
  _T_3_0_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _T_3_0_dirty = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_3_1_tag = _RAND_4[16:0];
  _RAND_5 = {1{`RANDOM}};
  _T_3_1_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _T_3_1_dirty = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_3_2_tag = _RAND_7[16:0];
  _RAND_8 = {1{`RANDOM}};
  _T_3_2_valid = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _T_3_2_dirty = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _T_3_3_tag = _RAND_10[16:0];
  _RAND_11 = {1{`RANDOM}};
  _T_3_3_valid = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _T_3_3_dirty = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_1 <= io_r_0_req_ready & io_r_0_req_valid;
    if (reset) begin
      _T_3_0_tag <= 17'h0;
    end else if (_T_1) begin
      _T_3_0_tag <= ram_io_r_resp_data_0_tag;
    end
    if (reset) begin
      _T_3_0_valid <= 1'h0;
    end else if (_T_1) begin
      _T_3_0_valid <= ram_io_r_resp_data_0_valid;
    end
    if (reset) begin
      _T_3_0_dirty <= 1'h0;
    end else if (_T_1) begin
      _T_3_0_dirty <= ram_io_r_resp_data_0_dirty;
    end
    if (reset) begin
      _T_3_1_tag <= 17'h0;
    end else if (_T_1) begin
      _T_3_1_tag <= ram_io_r_resp_data_1_tag;
    end
    if (reset) begin
      _T_3_1_valid <= 1'h0;
    end else if (_T_1) begin
      _T_3_1_valid <= ram_io_r_resp_data_1_valid;
    end
    if (reset) begin
      _T_3_1_dirty <= 1'h0;
    end else if (_T_1) begin
      _T_3_1_dirty <= ram_io_r_resp_data_1_dirty;
    end
    if (reset) begin
      _T_3_2_tag <= 17'h0;
    end else if (_T_1) begin
      _T_3_2_tag <= ram_io_r_resp_data_2_tag;
    end
    if (reset) begin
      _T_3_2_valid <= 1'h0;
    end else if (_T_1) begin
      _T_3_2_valid <= ram_io_r_resp_data_2_valid;
    end
    if (reset) begin
      _T_3_2_dirty <= 1'h0;
    end else if (_T_1) begin
      _T_3_2_dirty <= ram_io_r_resp_data_2_dirty;
    end
    if (reset) begin
      _T_3_3_tag <= 17'h0;
    end else if (_T_1) begin
      _T_3_3_tag <= ram_io_r_resp_data_3_tag;
    end
    if (reset) begin
      _T_3_3_valid <= 1'h0;
    end else if (_T_1) begin
      _T_3_3_valid <= ram_io_r_resp_data_3_valid;
    end
    if (reset) begin
      _T_3_3_dirty <= 1'h0;
    end else if (_T_1) begin
      _T_3_3_dirty <= ram_io_r_resp_data_3_dirty;
    end
  end
endmodule
module SRAMTemplate_6(
  input         clock,
  output        io_r_req_ready,
  input         io_r_req_valid,
  input  [11:0] io_r_req_bits_setIdx,
  output [63:0] io_r_resp_data_0_data,
  output [63:0] io_r_resp_data_1_data,
  output [63:0] io_r_resp_data_2_data,
  output [63:0] io_r_resp_data_3_data,
  input         io_w_req_valid,
  input  [11:0] io_w_req_bits_setIdx,
  input  [63:0] io_w_req_bits_data_data,
  input  [3:0]  io_w_req_bits_waymask
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_9;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] array_0 [0:4095]; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_0__T_13_data; // @[SRAMTemplate.scala 76:26]
  wire [11:0] array_0__T_13_addr; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_0__T_9_data; // @[SRAMTemplate.scala 76:26]
  wire [11:0] array_0__T_9_addr; // @[SRAMTemplate.scala 76:26]
  wire  array_0__T_9_mask; // @[SRAMTemplate.scala 76:26]
  wire  array_0__T_9_en; // @[SRAMTemplate.scala 76:26]
  reg  array_0__T_13_en_pipe_0;
  reg [11:0] array_0__T_13_addr_pipe_0;
  reg [63:0] array_1 [0:4095]; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_1__T_13_data; // @[SRAMTemplate.scala 76:26]
  wire [11:0] array_1__T_13_addr; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_1__T_9_data; // @[SRAMTemplate.scala 76:26]
  wire [11:0] array_1__T_9_addr; // @[SRAMTemplate.scala 76:26]
  wire  array_1__T_9_mask; // @[SRAMTemplate.scala 76:26]
  wire  array_1__T_9_en; // @[SRAMTemplate.scala 76:26]
  reg  array_1__T_13_en_pipe_0;
  reg [11:0] array_1__T_13_addr_pipe_0;
  reg [63:0] array_2 [0:4095]; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_2__T_13_data; // @[SRAMTemplate.scala 76:26]
  wire [11:0] array_2__T_13_addr; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_2__T_9_data; // @[SRAMTemplate.scala 76:26]
  wire [11:0] array_2__T_9_addr; // @[SRAMTemplate.scala 76:26]
  wire  array_2__T_9_mask; // @[SRAMTemplate.scala 76:26]
  wire  array_2__T_9_en; // @[SRAMTemplate.scala 76:26]
  reg  array_2__T_13_en_pipe_0;
  reg [11:0] array_2__T_13_addr_pipe_0;
  reg [63:0] array_3 [0:4095]; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_3__T_13_data; // @[SRAMTemplate.scala 76:26]
  wire [11:0] array_3__T_13_addr; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_3__T_9_data; // @[SRAMTemplate.scala 76:26]
  wire [11:0] array_3__T_9_addr; // @[SRAMTemplate.scala 76:26]
  wire  array_3__T_9_mask; // @[SRAMTemplate.scala 76:26]
  wire  array_3__T_9_en; // @[SRAMTemplate.scala 76:26]
  reg  array_3__T_13_en_pipe_0;
  reg [11:0] array_3__T_13_addr_pipe_0;
  wire  _T = ~io_w_req_valid; // @[SRAMTemplate.scala 89:41]
  assign array_0__T_13_addr = array_0__T_13_addr_pipe_0;
  assign array_0__T_13_data = array_0[array_0__T_13_addr]; // @[SRAMTemplate.scala 76:26]
  assign array_0__T_9_data = io_w_req_bits_data_data;
  assign array_0__T_9_addr = io_w_req_bits_setIdx;
  assign array_0__T_9_mask = io_w_req_bits_waymask[0];
  assign array_0__T_9_en = io_w_req_valid;
  assign array_1__T_13_addr = array_1__T_13_addr_pipe_0;
  assign array_1__T_13_data = array_1[array_1__T_13_addr]; // @[SRAMTemplate.scala 76:26]
  assign array_1__T_9_data = io_w_req_bits_data_data;
  assign array_1__T_9_addr = io_w_req_bits_setIdx;
  assign array_1__T_9_mask = io_w_req_bits_waymask[1];
  assign array_1__T_9_en = io_w_req_valid;
  assign array_2__T_13_addr = array_2__T_13_addr_pipe_0;
  assign array_2__T_13_data = array_2[array_2__T_13_addr]; // @[SRAMTemplate.scala 76:26]
  assign array_2__T_9_data = io_w_req_bits_data_data;
  assign array_2__T_9_addr = io_w_req_bits_setIdx;
  assign array_2__T_9_mask = io_w_req_bits_waymask[2];
  assign array_2__T_9_en = io_w_req_valid;
  assign array_3__T_13_addr = array_3__T_13_addr_pipe_0;
  assign array_3__T_13_data = array_3[array_3__T_13_addr]; // @[SRAMTemplate.scala 76:26]
  assign array_3__T_9_data = io_w_req_bits_data_data;
  assign array_3__T_9_addr = io_w_req_bits_setIdx;
  assign array_3__T_9_mask = io_w_req_bits_waymask[3];
  assign array_3__T_9_en = io_w_req_valid;
  assign io_r_req_ready = ~io_w_req_valid; // @[SRAMTemplate.scala 101:18]
  assign io_r_resp_data_0_data = array_0__T_13_data; // @[SRAMTemplate.scala 99:18]
  assign io_r_resp_data_1_data = array_1__T_13_data; // @[SRAMTemplate.scala 99:18]
  assign io_r_resp_data_2_data = array_2__T_13_data; // @[SRAMTemplate.scala 99:18]
  assign io_r_resp_data_3_data = array_3__T_13_data; // @[SRAMTemplate.scala 99:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4096; initvar = initvar+1)
    array_0[initvar] = _RAND_0[63:0];
  _RAND_3 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4096; initvar = initvar+1)
    array_1[initvar] = _RAND_3[63:0];
  _RAND_6 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4096; initvar = initvar+1)
    array_2[initvar] = _RAND_6[63:0];
  _RAND_9 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4096; initvar = initvar+1)
    array_3[initvar] = _RAND_9[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  array_0__T_13_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  array_0__T_13_addr_pipe_0 = _RAND_2[11:0];
  _RAND_4 = {1{`RANDOM}};
  array_1__T_13_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  array_1__T_13_addr_pipe_0 = _RAND_5[11:0];
  _RAND_7 = {1{`RANDOM}};
  array_2__T_13_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  array_2__T_13_addr_pipe_0 = _RAND_8[11:0];
  _RAND_10 = {1{`RANDOM}};
  array_3__T_13_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  array_3__T_13_addr_pipe_0 = _RAND_11[11:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(array_0__T_9_en & array_0__T_9_mask) begin
      array_0[array_0__T_9_addr] <= array_0__T_9_data; // @[SRAMTemplate.scala 76:26]
    end
    array_0__T_13_en_pipe_0 <= io_r_req_valid & _T;
    if (io_r_req_valid & _T) begin
      array_0__T_13_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if(array_1__T_9_en & array_1__T_9_mask) begin
      array_1[array_1__T_9_addr] <= array_1__T_9_data; // @[SRAMTemplate.scala 76:26]
    end
    array_1__T_13_en_pipe_0 <= io_r_req_valid & _T;
    if (io_r_req_valid & _T) begin
      array_1__T_13_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if(array_2__T_9_en & array_2__T_9_mask) begin
      array_2[array_2__T_9_addr] <= array_2__T_9_data; // @[SRAMTemplate.scala 76:26]
    end
    array_2__T_13_en_pipe_0 <= io_r_req_valid & _T;
    if (io_r_req_valid & _T) begin
      array_2__T_13_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
    if(array_3__T_9_en & array_3__T_9_mask) begin
      array_3[array_3__T_9_addr] <= array_3__T_9_data; // @[SRAMTemplate.scala 76:26]
    end
    array_3__T_13_en_pipe_0 <= io_r_req_valid & _T;
    if (io_r_req_valid & _T) begin
      array_3__T_13_addr_pipe_0 <= io_r_req_bits_setIdx;
    end
  end
endmodule
module Arbiter_13(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [11:0] io_in_0_bits_setIdx,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [11:0] io_in_1_bits_setIdx,
  input         io_out_ready,
  output        io_out_valid,
  output [11:0] io_out_bits_setIdx
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  wire  _T_2 = ~grant_1; // @[Arbiter.scala 135:19]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:14]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_out_valid = _T_2 | io_in_1_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
endmodule
module SRAMTemplateWithArbiter_5(
  input         clock,
  input         reset,
  output        io_r_0_req_ready,
  input         io_r_0_req_valid,
  input  [11:0] io_r_0_req_bits_setIdx,
  output [63:0] io_r_0_resp_data_0_data,
  output [63:0] io_r_0_resp_data_1_data,
  output [63:0] io_r_0_resp_data_2_data,
  output [63:0] io_r_0_resp_data_3_data,
  output        io_r_1_req_ready,
  input         io_r_1_req_valid,
  input  [11:0] io_r_1_req_bits_setIdx,
  output [63:0] io_r_1_resp_data_0_data,
  output [63:0] io_r_1_resp_data_1_data,
  output [63:0] io_r_1_resp_data_2_data,
  output [63:0] io_r_1_resp_data_3_data,
  input         io_w_req_valid,
  input  [11:0] io_w_req_bits_setIdx,
  input  [63:0] io_w_req_bits_data_data,
  input  [3:0]  io_w_req_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  ram_clock; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_r_req_ready; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_r_req_valid; // @[SRAMTemplate.scala 121:19]
  wire [11:0] ram_io_r_req_bits_setIdx; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_r_resp_data_0_data; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_r_resp_data_1_data; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_r_resp_data_2_data; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_r_resp_data_3_data; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_w_req_valid; // @[SRAMTemplate.scala 121:19]
  wire [11:0] ram_io_w_req_bits_setIdx; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_w_req_bits_data_data; // @[SRAMTemplate.scala 121:19]
  wire [3:0] ram_io_w_req_bits_waymask; // @[SRAMTemplate.scala 121:19]
  wire  readArb_io_in_0_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_in_0_valid; // @[SRAMTemplate.scala 124:23]
  wire [11:0] readArb_io_in_0_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_in_1_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_in_1_valid; // @[SRAMTemplate.scala 124:23]
  wire [11:0] readArb_io_in_1_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_out_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_out_valid; // @[SRAMTemplate.scala 124:23]
  wire [11:0] readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  reg  _T_1; // @[SRAMTemplate.scala 130:58]
  reg [63:0] _T_3_0_data; // @[Reg.scala 27:20]
  reg [63:0] _T_3_1_data; // @[Reg.scala 27:20]
  reg [63:0] _T_3_2_data; // @[Reg.scala 27:20]
  reg [63:0] _T_3_3_data; // @[Reg.scala 27:20]
  reg  _T_6; // @[SRAMTemplate.scala 130:58]
  reg [63:0] _T_8_0_data; // @[Reg.scala 27:20]
  reg [63:0] _T_8_1_data; // @[Reg.scala 27:20]
  reg [63:0] _T_8_2_data; // @[Reg.scala 27:20]
  reg [63:0] _T_8_3_data; // @[Reg.scala 27:20]
  SRAMTemplate_6 ram ( // @[SRAMTemplate.scala 121:19]
    .clock(ram_clock),
    .io_r_req_ready(ram_io_r_req_ready),
    .io_r_req_valid(ram_io_r_req_valid),
    .io_r_req_bits_setIdx(ram_io_r_req_bits_setIdx),
    .io_r_resp_data_0_data(ram_io_r_resp_data_0_data),
    .io_r_resp_data_1_data(ram_io_r_resp_data_1_data),
    .io_r_resp_data_2_data(ram_io_r_resp_data_2_data),
    .io_r_resp_data_3_data(ram_io_r_resp_data_3_data),
    .io_w_req_valid(ram_io_w_req_valid),
    .io_w_req_bits_setIdx(ram_io_w_req_bits_setIdx),
    .io_w_req_bits_data_data(ram_io_w_req_bits_data_data),
    .io_w_req_bits_waymask(ram_io_w_req_bits_waymask)
  );
  Arbiter_13 readArb ( // @[SRAMTemplate.scala 124:23]
    .io_in_0_ready(readArb_io_in_0_ready),
    .io_in_0_valid(readArb_io_in_0_valid),
    .io_in_0_bits_setIdx(readArb_io_in_0_bits_setIdx),
    .io_in_1_ready(readArb_io_in_1_ready),
    .io_in_1_valid(readArb_io_in_1_valid),
    .io_in_1_bits_setIdx(readArb_io_in_1_bits_setIdx),
    .io_out_ready(readArb_io_out_ready),
    .io_out_valid(readArb_io_out_valid),
    .io_out_bits_setIdx(readArb_io_out_bits_setIdx)
  );
  assign io_r_0_req_ready = readArb_io_in_0_ready; // @[SRAMTemplate.scala 125:17]
  assign io_r_0_resp_data_0_data = _T_1 ? ram_io_r_resp_data_0_data : _T_3_0_data; // @[SRAMTemplate.scala 130:17]
  assign io_r_0_resp_data_1_data = _T_1 ? ram_io_r_resp_data_1_data : _T_3_1_data; // @[SRAMTemplate.scala 130:17]
  assign io_r_0_resp_data_2_data = _T_1 ? ram_io_r_resp_data_2_data : _T_3_2_data; // @[SRAMTemplate.scala 130:17]
  assign io_r_0_resp_data_3_data = _T_1 ? ram_io_r_resp_data_3_data : _T_3_3_data; // @[SRAMTemplate.scala 130:17]
  assign io_r_1_req_ready = readArb_io_in_1_ready; // @[SRAMTemplate.scala 125:17]
  assign io_r_1_resp_data_0_data = _T_6 ? ram_io_r_resp_data_0_data : _T_8_0_data; // @[SRAMTemplate.scala 130:17]
  assign io_r_1_resp_data_1_data = _T_6 ? ram_io_r_resp_data_1_data : _T_8_1_data; // @[SRAMTemplate.scala 130:17]
  assign io_r_1_resp_data_2_data = _T_6 ? ram_io_r_resp_data_2_data : _T_8_2_data; // @[SRAMTemplate.scala 130:17]
  assign io_r_1_resp_data_3_data = _T_6 ? ram_io_r_resp_data_3_data : _T_8_3_data; // @[SRAMTemplate.scala 130:17]
  assign ram_clock = clock;
  assign ram_io_r_req_valid = readArb_io_out_valid; // @[SRAMTemplate.scala 126:16]
  assign ram_io_r_req_bits_setIdx = readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 126:16]
  assign ram_io_w_req_valid = io_w_req_valid; // @[SRAMTemplate.scala 122:12]
  assign ram_io_w_req_bits_setIdx = io_w_req_bits_setIdx; // @[SRAMTemplate.scala 122:12]
  assign ram_io_w_req_bits_data_data = io_w_req_bits_data_data; // @[SRAMTemplate.scala 122:12]
  assign ram_io_w_req_bits_waymask = io_w_req_bits_waymask; // @[SRAMTemplate.scala 122:12]
  assign readArb_io_in_0_valid = io_r_0_req_valid; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_in_0_bits_setIdx = io_r_0_req_bits_setIdx; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_in_1_valid = io_r_1_req_valid; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_in_1_bits_setIdx = io_r_1_req_bits_setIdx; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_out_ready = ram_io_r_req_ready; // @[SRAMTemplate.scala 126:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1 = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  _T_3_0_data = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  _T_3_1_data = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  _T_3_2_data = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  _T_3_3_data = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  _T_6 = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  _T_8_0_data = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  _T_8_1_data = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  _T_8_2_data = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  _T_8_3_data = _RAND_9[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_1 <= io_r_0_req_ready & io_r_0_req_valid;
    if (reset) begin
      _T_3_0_data <= 64'h0;
    end else if (_T_1) begin
      _T_3_0_data <= ram_io_r_resp_data_0_data;
    end
    if (reset) begin
      _T_3_1_data <= 64'h0;
    end else if (_T_1) begin
      _T_3_1_data <= ram_io_r_resp_data_1_data;
    end
    if (reset) begin
      _T_3_2_data <= 64'h0;
    end else if (_T_1) begin
      _T_3_2_data <= ram_io_r_resp_data_2_data;
    end
    if (reset) begin
      _T_3_3_data <= 64'h0;
    end else if (_T_1) begin
      _T_3_3_data <= ram_io_r_resp_data_3_data;
    end
    _T_6 <= io_r_1_req_ready & io_r_1_req_valid;
    if (reset) begin
      _T_8_0_data <= 64'h0;
    end else if (_T_6) begin
      _T_8_0_data <= ram_io_r_resp_data_0_data;
    end
    if (reset) begin
      _T_8_1_data <= 64'h0;
    end else if (_T_6) begin
      _T_8_1_data <= ram_io_r_resp_data_1_data;
    end
    if (reset) begin
      _T_8_2_data <= 64'h0;
    end else if (_T_6) begin
      _T_8_2_data <= ram_io_r_resp_data_2_data;
    end
    if (reset) begin
      _T_8_3_data <= 64'h0;
    end else if (_T_6) begin
      _T_8_3_data <= ram_io_r_resp_data_3_data;
    end
  end
endmodule
module Cache_2(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [2:0]  io_in_req_bits_size,
  input  [3:0]  io_in_req_bits_cmd,
  input  [7:0]  io_in_req_bits_wmask,
  input  [63:0] io_in_req_bits_wdata,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_mem_req_ready,
  output        io_out_mem_req_valid,
  output [31:0] io_out_mem_req_bits_addr,
  output [3:0]  io_out_mem_req_bits_cmd,
  output [63:0] io_out_mem_req_bits_wdata,
  input         io_out_mem_resp_valid,
  input  [3:0]  io_out_mem_resp_bits_cmd,
  input  [63:0] io_out_mem_resp_bits_rdata,
  input         DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
`endif // RANDOMIZE_REG_INIT
  wire  s1_clock; // @[Cache.scala 475:18]
  wire  s1_reset; // @[Cache.scala 475:18]
  wire  s1_io_in_ready; // @[Cache.scala 475:18]
  wire  s1_io_in_valid; // @[Cache.scala 475:18]
  wire [31:0] s1_io_in_bits_addr; // @[Cache.scala 475:18]
  wire [2:0] s1_io_in_bits_size; // @[Cache.scala 475:18]
  wire [3:0] s1_io_in_bits_cmd; // @[Cache.scala 475:18]
  wire [7:0] s1_io_in_bits_wmask; // @[Cache.scala 475:18]
  wire [63:0] s1_io_in_bits_wdata; // @[Cache.scala 475:18]
  wire  s1_io_out_ready; // @[Cache.scala 475:18]
  wire  s1_io_out_valid; // @[Cache.scala 475:18]
  wire [31:0] s1_io_out_bits_req_addr; // @[Cache.scala 475:18]
  wire [2:0] s1_io_out_bits_req_size; // @[Cache.scala 475:18]
  wire [3:0] s1_io_out_bits_req_cmd; // @[Cache.scala 475:18]
  wire [7:0] s1_io_out_bits_req_wmask; // @[Cache.scala 475:18]
  wire [63:0] s1_io_out_bits_req_wdata; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_req_ready; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_req_valid; // @[Cache.scala 475:18]
  wire [8:0] s1_io_metaReadBus_req_bits_setIdx; // @[Cache.scala 475:18]
  wire [16:0] s1_io_metaReadBus_resp_data_0_tag; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_0_valid; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_0_dirty; // @[Cache.scala 475:18]
  wire [16:0] s1_io_metaReadBus_resp_data_1_tag; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_1_valid; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_1_dirty; // @[Cache.scala 475:18]
  wire [16:0] s1_io_metaReadBus_resp_data_2_tag; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_2_valid; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_2_dirty; // @[Cache.scala 475:18]
  wire [16:0] s1_io_metaReadBus_resp_data_3_tag; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_3_valid; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_3_dirty; // @[Cache.scala 475:18]
  wire  s1_io_dataReadBus_req_ready; // @[Cache.scala 475:18]
  wire  s1_io_dataReadBus_req_valid; // @[Cache.scala 475:18]
  wire [11:0] s1_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 475:18]
  wire [63:0] s1_io_dataReadBus_resp_data_0_data; // @[Cache.scala 475:18]
  wire [63:0] s1_io_dataReadBus_resp_data_1_data; // @[Cache.scala 475:18]
  wire [63:0] s1_io_dataReadBus_resp_data_2_data; // @[Cache.scala 475:18]
  wire [63:0] s1_io_dataReadBus_resp_data_3_data; // @[Cache.scala 475:18]
  wire  s1_DISPLAY_ENABLE; // @[Cache.scala 475:18]
  wire  s2_clock; // @[Cache.scala 476:18]
  wire  s2_reset; // @[Cache.scala 476:18]
  wire  s2_io_in_ready; // @[Cache.scala 476:18]
  wire  s2_io_in_valid; // @[Cache.scala 476:18]
  wire [31:0] s2_io_in_bits_req_addr; // @[Cache.scala 476:18]
  wire [2:0] s2_io_in_bits_req_size; // @[Cache.scala 476:18]
  wire [3:0] s2_io_in_bits_req_cmd; // @[Cache.scala 476:18]
  wire [7:0] s2_io_in_bits_req_wmask; // @[Cache.scala 476:18]
  wire [63:0] s2_io_in_bits_req_wdata; // @[Cache.scala 476:18]
  wire  s2_io_out_ready; // @[Cache.scala 476:18]
  wire  s2_io_out_valid; // @[Cache.scala 476:18]
  wire [31:0] s2_io_out_bits_req_addr; // @[Cache.scala 476:18]
  wire [2:0] s2_io_out_bits_req_size; // @[Cache.scala 476:18]
  wire [3:0] s2_io_out_bits_req_cmd; // @[Cache.scala 476:18]
  wire [7:0] s2_io_out_bits_req_wmask; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_req_wdata; // @[Cache.scala 476:18]
  wire [16:0] s2_io_out_bits_metas_0_tag; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_0_valid; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_0_dirty; // @[Cache.scala 476:18]
  wire [16:0] s2_io_out_bits_metas_1_tag; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_1_valid; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_1_dirty; // @[Cache.scala 476:18]
  wire [16:0] s2_io_out_bits_metas_2_tag; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_2_valid; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_2_dirty; // @[Cache.scala 476:18]
  wire [16:0] s2_io_out_bits_metas_3_tag; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_3_valid; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_3_dirty; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_datas_0_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_datas_1_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_datas_2_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_datas_3_data; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_hit; // @[Cache.scala 476:18]
  wire [3:0] s2_io_out_bits_waymask; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_mmio; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_isForwardData; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_forwardData_data_data; // @[Cache.scala 476:18]
  wire [3:0] s2_io_out_bits_forwardData_waymask; // @[Cache.scala 476:18]
  wire [16:0] s2_io_metaReadResp_0_tag; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_0_valid; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_0_dirty; // @[Cache.scala 476:18]
  wire [16:0] s2_io_metaReadResp_1_tag; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_1_valid; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_1_dirty; // @[Cache.scala 476:18]
  wire [16:0] s2_io_metaReadResp_2_tag; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_2_valid; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_2_dirty; // @[Cache.scala 476:18]
  wire [16:0] s2_io_metaReadResp_3_tag; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_3_valid; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_3_dirty; // @[Cache.scala 476:18]
  wire [63:0] s2_io_dataReadResp_0_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_dataReadResp_1_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_dataReadResp_2_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_dataReadResp_3_data; // @[Cache.scala 476:18]
  wire  s2_io_metaWriteBus_req_valid; // @[Cache.scala 476:18]
  wire [8:0] s2_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 476:18]
  wire [16:0] s2_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 476:18]
  wire  s2_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 476:18]
  wire [3:0] s2_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 476:18]
  wire  s2_io_dataWriteBus_req_valid; // @[Cache.scala 476:18]
  wire [11:0] s2_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 476:18]
  wire [63:0] s2_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 476:18]
  wire [3:0] s2_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 476:18]
  wire  s2_DISPLAY_ENABLE; // @[Cache.scala 476:18]
  wire  s3_clock; // @[Cache.scala 477:18]
  wire  s3_reset; // @[Cache.scala 477:18]
  wire  s3_io_in_ready; // @[Cache.scala 477:18]
  wire  s3_io_in_valid; // @[Cache.scala 477:18]
  wire [31:0] s3_io_in_bits_req_addr; // @[Cache.scala 477:18]
  wire [2:0] s3_io_in_bits_req_size; // @[Cache.scala 477:18]
  wire [3:0] s3_io_in_bits_req_cmd; // @[Cache.scala 477:18]
  wire [7:0] s3_io_in_bits_req_wmask; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_req_wdata; // @[Cache.scala 477:18]
  wire [16:0] s3_io_in_bits_metas_0_tag; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_0_valid; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_0_dirty; // @[Cache.scala 477:18]
  wire [16:0] s3_io_in_bits_metas_1_tag; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_1_valid; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_1_dirty; // @[Cache.scala 477:18]
  wire [16:0] s3_io_in_bits_metas_2_tag; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_2_valid; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_2_dirty; // @[Cache.scala 477:18]
  wire [16:0] s3_io_in_bits_metas_3_tag; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_3_valid; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_3_dirty; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_datas_0_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_datas_1_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_datas_2_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_datas_3_data; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_hit; // @[Cache.scala 477:18]
  wire [3:0] s3_io_in_bits_waymask; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_mmio; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_isForwardData; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_forwardData_data_data; // @[Cache.scala 477:18]
  wire [3:0] s3_io_in_bits_forwardData_waymask; // @[Cache.scala 477:18]
  wire  s3_io_out_ready; // @[Cache.scala 477:18]
  wire  s3_io_out_valid; // @[Cache.scala 477:18]
  wire [3:0] s3_io_out_bits_cmd; // @[Cache.scala 477:18]
  wire [63:0] s3_io_out_bits_rdata; // @[Cache.scala 477:18]
  wire  s3_io_isFinish; // @[Cache.scala 477:18]
  wire  s3_io_dataReadBus_req_ready; // @[Cache.scala 477:18]
  wire  s3_io_dataReadBus_req_valid; // @[Cache.scala 477:18]
  wire [11:0] s3_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 477:18]
  wire [63:0] s3_io_dataReadBus_resp_data_0_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_dataReadBus_resp_data_1_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_dataReadBus_resp_data_2_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_dataReadBus_resp_data_3_data; // @[Cache.scala 477:18]
  wire  s3_io_dataWriteBus_req_valid; // @[Cache.scala 477:18]
  wire [11:0] s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 477:18]
  wire [63:0] s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 477:18]
  wire [3:0] s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 477:18]
  wire  s3_io_metaWriteBus_req_valid; // @[Cache.scala 477:18]
  wire [8:0] s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 477:18]
  wire [16:0] s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 477:18]
  wire  s3_io_metaWriteBus_req_bits_data_valid; // @[Cache.scala 477:18]
  wire  s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 477:18]
  wire [3:0] s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 477:18]
  wire  s3_io_mem_req_ready; // @[Cache.scala 477:18]
  wire  s3_io_mem_req_valid; // @[Cache.scala 477:18]
  wire [31:0] s3_io_mem_req_bits_addr; // @[Cache.scala 477:18]
  wire [2:0] s3_io_mem_req_bits_size; // @[Cache.scala 477:18]
  wire [3:0] s3_io_mem_req_bits_cmd; // @[Cache.scala 477:18]
  wire [7:0] s3_io_mem_req_bits_wmask; // @[Cache.scala 477:18]
  wire [63:0] s3_io_mem_req_bits_wdata; // @[Cache.scala 477:18]
  wire  s3_io_mem_resp_ready; // @[Cache.scala 477:18]
  wire  s3_io_mem_resp_valid; // @[Cache.scala 477:18]
  wire [3:0] s3_io_mem_resp_bits_cmd; // @[Cache.scala 477:18]
  wire [63:0] s3_io_mem_resp_bits_rdata; // @[Cache.scala 477:18]
  wire  s3_io_cohResp_valid; // @[Cache.scala 477:18]
  wire  s3_io_dataReadRespToL1; // @[Cache.scala 477:18]
  wire  s3_DISPLAY_ENABLE; // @[Cache.scala 477:18]
  wire  metaArray_clock; // @[Cache.scala 478:25]
  wire  metaArray_reset; // @[Cache.scala 478:25]
  wire  metaArray_io_r_0_req_ready; // @[Cache.scala 478:25]
  wire  metaArray_io_r_0_req_valid; // @[Cache.scala 478:25]
  wire [8:0] metaArray_io_r_0_req_bits_setIdx; // @[Cache.scala 478:25]
  wire [16:0] metaArray_io_r_0_resp_data_0_tag; // @[Cache.scala 478:25]
  wire  metaArray_io_r_0_resp_data_0_valid; // @[Cache.scala 478:25]
  wire  metaArray_io_r_0_resp_data_0_dirty; // @[Cache.scala 478:25]
  wire [16:0] metaArray_io_r_0_resp_data_1_tag; // @[Cache.scala 478:25]
  wire  metaArray_io_r_0_resp_data_1_valid; // @[Cache.scala 478:25]
  wire  metaArray_io_r_0_resp_data_1_dirty; // @[Cache.scala 478:25]
  wire [16:0] metaArray_io_r_0_resp_data_2_tag; // @[Cache.scala 478:25]
  wire  metaArray_io_r_0_resp_data_2_valid; // @[Cache.scala 478:25]
  wire  metaArray_io_r_0_resp_data_2_dirty; // @[Cache.scala 478:25]
  wire [16:0] metaArray_io_r_0_resp_data_3_tag; // @[Cache.scala 478:25]
  wire  metaArray_io_r_0_resp_data_3_valid; // @[Cache.scala 478:25]
  wire  metaArray_io_r_0_resp_data_3_dirty; // @[Cache.scala 478:25]
  wire  metaArray_io_w_req_valid; // @[Cache.scala 478:25]
  wire [8:0] metaArray_io_w_req_bits_setIdx; // @[Cache.scala 478:25]
  wire [16:0] metaArray_io_w_req_bits_data_tag; // @[Cache.scala 478:25]
  wire  metaArray_io_w_req_bits_data_dirty; // @[Cache.scala 478:25]
  wire [3:0] metaArray_io_w_req_bits_waymask; // @[Cache.scala 478:25]
  wire  dataArray_clock; // @[Cache.scala 479:25]
  wire  dataArray_reset; // @[Cache.scala 479:25]
  wire  dataArray_io_r_0_req_ready; // @[Cache.scala 479:25]
  wire  dataArray_io_r_0_req_valid; // @[Cache.scala 479:25]
  wire [11:0] dataArray_io_r_0_req_bits_setIdx; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r_0_resp_data_0_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r_0_resp_data_1_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r_0_resp_data_2_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r_0_resp_data_3_data; // @[Cache.scala 479:25]
  wire  dataArray_io_r_1_req_ready; // @[Cache.scala 479:25]
  wire  dataArray_io_r_1_req_valid; // @[Cache.scala 479:25]
  wire [11:0] dataArray_io_r_1_req_bits_setIdx; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r_1_resp_data_0_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r_1_resp_data_1_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r_1_resp_data_2_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r_1_resp_data_3_data; // @[Cache.scala 479:25]
  wire  dataArray_io_w_req_valid; // @[Cache.scala 479:25]
  wire [11:0] dataArray_io_w_req_bits_setIdx; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_w_req_bits_data_data; // @[Cache.scala 479:25]
  wire [3:0] dataArray_io_w_req_bits_waymask; // @[Cache.scala 479:25]
  wire  arb_io_in_0_ready; // @[Cache.scala 488:19]
  wire  arb_io_in_0_valid; // @[Cache.scala 488:19]
  wire [31:0] arb_io_in_0_bits_addr; // @[Cache.scala 488:19]
  wire [2:0] arb_io_in_0_bits_size; // @[Cache.scala 488:19]
  wire [3:0] arb_io_in_0_bits_cmd; // @[Cache.scala 488:19]
  wire [7:0] arb_io_in_0_bits_wmask; // @[Cache.scala 488:19]
  wire [63:0] arb_io_in_0_bits_wdata; // @[Cache.scala 488:19]
  wire  arb_io_in_1_ready; // @[Cache.scala 488:19]
  wire  arb_io_in_1_valid; // @[Cache.scala 488:19]
  wire [31:0] arb_io_in_1_bits_addr; // @[Cache.scala 488:19]
  wire [2:0] arb_io_in_1_bits_size; // @[Cache.scala 488:19]
  wire [3:0] arb_io_in_1_bits_cmd; // @[Cache.scala 488:19]
  wire [7:0] arb_io_in_1_bits_wmask; // @[Cache.scala 488:19]
  wire [63:0] arb_io_in_1_bits_wdata; // @[Cache.scala 488:19]
  wire  arb_io_out_ready; // @[Cache.scala 488:19]
  wire  arb_io_out_valid; // @[Cache.scala 488:19]
  wire [31:0] arb_io_out_bits_addr; // @[Cache.scala 488:19]
  wire [2:0] arb_io_out_bits_size; // @[Cache.scala 488:19]
  wire [3:0] arb_io_out_bits_cmd; // @[Cache.scala 488:19]
  wire [7:0] arb_io_out_bits_wmask; // @[Cache.scala 488:19]
  wire [63:0] arb_io_out_bits_wdata; // @[Cache.scala 488:19]
  wire  _T = s2_io_out_ready & s2_io_out_valid; // @[Decoupled.scala 40:37]
  reg  _T_2; // @[Pipeline.scala 24:24]
  wire  _GEN_0 = _T ? 1'h0 : _T_2; // @[Pipeline.scala 25:25]
  wire  _T_3 = s1_io_out_valid & s2_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_1 = _T_3 | _GEN_0; // @[Pipeline.scala 26:38]
  reg [31:0] _T_5_req_addr; // @[Reg.scala 15:16]
  reg [2:0] _T_5_req_size; // @[Reg.scala 15:16]
  reg [3:0] _T_5_req_cmd; // @[Reg.scala 15:16]
  reg [7:0] _T_5_req_wmask; // @[Reg.scala 15:16]
  reg [63:0] _T_5_req_wdata; // @[Reg.scala 15:16]
  reg  _T_7; // @[Pipeline.scala 24:24]
  wire  _GEN_8 = s3_io_isFinish ? 1'h0 : _T_7; // @[Pipeline.scala 25:25]
  wire  _T_8 = s2_io_out_valid & s3_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_9 = _T_8 | _GEN_8; // @[Pipeline.scala 26:38]
  reg [31:0] _T_10_req_addr; // @[Reg.scala 15:16]
  reg [2:0] _T_10_req_size; // @[Reg.scala 15:16]
  reg [3:0] _T_10_req_cmd; // @[Reg.scala 15:16]
  reg [7:0] _T_10_req_wmask; // @[Reg.scala 15:16]
  reg [63:0] _T_10_req_wdata; // @[Reg.scala 15:16]
  reg [16:0] _T_10_metas_0_tag; // @[Reg.scala 15:16]
  reg  _T_10_metas_0_valid; // @[Reg.scala 15:16]
  reg  _T_10_metas_0_dirty; // @[Reg.scala 15:16]
  reg [16:0] _T_10_metas_1_tag; // @[Reg.scala 15:16]
  reg  _T_10_metas_1_valid; // @[Reg.scala 15:16]
  reg  _T_10_metas_1_dirty; // @[Reg.scala 15:16]
  reg [16:0] _T_10_metas_2_tag; // @[Reg.scala 15:16]
  reg  _T_10_metas_2_valid; // @[Reg.scala 15:16]
  reg  _T_10_metas_2_dirty; // @[Reg.scala 15:16]
  reg [16:0] _T_10_metas_3_tag; // @[Reg.scala 15:16]
  reg  _T_10_metas_3_valid; // @[Reg.scala 15:16]
  reg  _T_10_metas_3_dirty; // @[Reg.scala 15:16]
  reg [63:0] _T_10_datas_0_data; // @[Reg.scala 15:16]
  reg [63:0] _T_10_datas_1_data; // @[Reg.scala 15:16]
  reg [63:0] _T_10_datas_2_data; // @[Reg.scala 15:16]
  reg [63:0] _T_10_datas_3_data; // @[Reg.scala 15:16]
  reg  _T_10_hit; // @[Reg.scala 15:16]
  reg [3:0] _T_10_waymask; // @[Reg.scala 15:16]
  reg  _T_10_mmio; // @[Reg.scala 15:16]
  reg  _T_10_isForwardData; // @[Reg.scala 15:16]
  reg [63:0] _T_10_forwardData_data_data; // @[Reg.scala 15:16]
  reg [3:0] _T_10_forwardData_waymask; // @[Reg.scala 15:16]
  wire  _T_15 = s3_io_out_bits_cmd == 4'h4; // @[SimpleBus.scala 95:26]
  wire  _T_16 = s3_io_out_valid & _T_15; // @[Cache.scala 505:43]
  wire  _T_17 = s3_io_out_valid | s3_io_dataReadRespToL1; // @[Cache.scala 505:100]
  reg [63:0] _T_20; // @[GTimer.scala 24:20]
  wire [63:0] _T_22 = _T_20 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_26 = ~reset; // @[Debug.scala 56:24]
  reg [63:0] _T_29; // @[GTimer.scala 24:20]
  wire [63:0] _T_31 = _T_29 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_38; // @[GTimer.scala 24:20]
  wire [63:0] _T_40 = _T_38 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_47; // @[GTimer.scala 24:20]
  wire [63:0] _T_49 = _T_47 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_56; // @[GTimer.scala 24:20]
  wire [63:0] _T_58 = _T_56 + 64'h1; // @[GTimer.scala 25:12]
  wire  _GEN_39 = s1_io_in_valid & DISPLAY_ENABLE; // @[Debug.scala 56:24]
  wire  _GEN_41 = s2_io_in_valid & DISPLAY_ENABLE; // @[Debug.scala 56:24]
  wire  _GEN_43 = s3_io_in_valid & DISPLAY_ENABLE; // @[Debug.scala 56:24]
  CacheStage1_2 s1 ( // @[Cache.scala 475:18]
    .clock(s1_clock),
    .reset(s1_reset),
    .io_in_ready(s1_io_in_ready),
    .io_in_valid(s1_io_in_valid),
    .io_in_bits_addr(s1_io_in_bits_addr),
    .io_in_bits_size(s1_io_in_bits_size),
    .io_in_bits_cmd(s1_io_in_bits_cmd),
    .io_in_bits_wmask(s1_io_in_bits_wmask),
    .io_in_bits_wdata(s1_io_in_bits_wdata),
    .io_out_ready(s1_io_out_ready),
    .io_out_valid(s1_io_out_valid),
    .io_out_bits_req_addr(s1_io_out_bits_req_addr),
    .io_out_bits_req_size(s1_io_out_bits_req_size),
    .io_out_bits_req_cmd(s1_io_out_bits_req_cmd),
    .io_out_bits_req_wmask(s1_io_out_bits_req_wmask),
    .io_out_bits_req_wdata(s1_io_out_bits_req_wdata),
    .io_metaReadBus_req_ready(s1_io_metaReadBus_req_ready),
    .io_metaReadBus_req_valid(s1_io_metaReadBus_req_valid),
    .io_metaReadBus_req_bits_setIdx(s1_io_metaReadBus_req_bits_setIdx),
    .io_metaReadBus_resp_data_0_tag(s1_io_metaReadBus_resp_data_0_tag),
    .io_metaReadBus_resp_data_0_valid(s1_io_metaReadBus_resp_data_0_valid),
    .io_metaReadBus_resp_data_0_dirty(s1_io_metaReadBus_resp_data_0_dirty),
    .io_metaReadBus_resp_data_1_tag(s1_io_metaReadBus_resp_data_1_tag),
    .io_metaReadBus_resp_data_1_valid(s1_io_metaReadBus_resp_data_1_valid),
    .io_metaReadBus_resp_data_1_dirty(s1_io_metaReadBus_resp_data_1_dirty),
    .io_metaReadBus_resp_data_2_tag(s1_io_metaReadBus_resp_data_2_tag),
    .io_metaReadBus_resp_data_2_valid(s1_io_metaReadBus_resp_data_2_valid),
    .io_metaReadBus_resp_data_2_dirty(s1_io_metaReadBus_resp_data_2_dirty),
    .io_metaReadBus_resp_data_3_tag(s1_io_metaReadBus_resp_data_3_tag),
    .io_metaReadBus_resp_data_3_valid(s1_io_metaReadBus_resp_data_3_valid),
    .io_metaReadBus_resp_data_3_dirty(s1_io_metaReadBus_resp_data_3_dirty),
    .io_dataReadBus_req_ready(s1_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s1_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s1_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s1_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s1_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s1_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s1_io_dataReadBus_resp_data_3_data),
    .DISPLAY_ENABLE(s1_DISPLAY_ENABLE)
  );
  CacheStage2_2 s2 ( // @[Cache.scala 476:18]
    .clock(s2_clock),
    .reset(s2_reset),
    .io_in_ready(s2_io_in_ready),
    .io_in_valid(s2_io_in_valid),
    .io_in_bits_req_addr(s2_io_in_bits_req_addr),
    .io_in_bits_req_size(s2_io_in_bits_req_size),
    .io_in_bits_req_cmd(s2_io_in_bits_req_cmd),
    .io_in_bits_req_wmask(s2_io_in_bits_req_wmask),
    .io_in_bits_req_wdata(s2_io_in_bits_req_wdata),
    .io_out_ready(s2_io_out_ready),
    .io_out_valid(s2_io_out_valid),
    .io_out_bits_req_addr(s2_io_out_bits_req_addr),
    .io_out_bits_req_size(s2_io_out_bits_req_size),
    .io_out_bits_req_cmd(s2_io_out_bits_req_cmd),
    .io_out_bits_req_wmask(s2_io_out_bits_req_wmask),
    .io_out_bits_req_wdata(s2_io_out_bits_req_wdata),
    .io_out_bits_metas_0_tag(s2_io_out_bits_metas_0_tag),
    .io_out_bits_metas_0_valid(s2_io_out_bits_metas_0_valid),
    .io_out_bits_metas_0_dirty(s2_io_out_bits_metas_0_dirty),
    .io_out_bits_metas_1_tag(s2_io_out_bits_metas_1_tag),
    .io_out_bits_metas_1_valid(s2_io_out_bits_metas_1_valid),
    .io_out_bits_metas_1_dirty(s2_io_out_bits_metas_1_dirty),
    .io_out_bits_metas_2_tag(s2_io_out_bits_metas_2_tag),
    .io_out_bits_metas_2_valid(s2_io_out_bits_metas_2_valid),
    .io_out_bits_metas_2_dirty(s2_io_out_bits_metas_2_dirty),
    .io_out_bits_metas_3_tag(s2_io_out_bits_metas_3_tag),
    .io_out_bits_metas_3_valid(s2_io_out_bits_metas_3_valid),
    .io_out_bits_metas_3_dirty(s2_io_out_bits_metas_3_dirty),
    .io_out_bits_datas_0_data(s2_io_out_bits_datas_0_data),
    .io_out_bits_datas_1_data(s2_io_out_bits_datas_1_data),
    .io_out_bits_datas_2_data(s2_io_out_bits_datas_2_data),
    .io_out_bits_datas_3_data(s2_io_out_bits_datas_3_data),
    .io_out_bits_hit(s2_io_out_bits_hit),
    .io_out_bits_waymask(s2_io_out_bits_waymask),
    .io_out_bits_mmio(s2_io_out_bits_mmio),
    .io_out_bits_isForwardData(s2_io_out_bits_isForwardData),
    .io_out_bits_forwardData_data_data(s2_io_out_bits_forwardData_data_data),
    .io_out_bits_forwardData_waymask(s2_io_out_bits_forwardData_waymask),
    .io_metaReadResp_0_tag(s2_io_metaReadResp_0_tag),
    .io_metaReadResp_0_valid(s2_io_metaReadResp_0_valid),
    .io_metaReadResp_0_dirty(s2_io_metaReadResp_0_dirty),
    .io_metaReadResp_1_tag(s2_io_metaReadResp_1_tag),
    .io_metaReadResp_1_valid(s2_io_metaReadResp_1_valid),
    .io_metaReadResp_1_dirty(s2_io_metaReadResp_1_dirty),
    .io_metaReadResp_2_tag(s2_io_metaReadResp_2_tag),
    .io_metaReadResp_2_valid(s2_io_metaReadResp_2_valid),
    .io_metaReadResp_2_dirty(s2_io_metaReadResp_2_dirty),
    .io_metaReadResp_3_tag(s2_io_metaReadResp_3_tag),
    .io_metaReadResp_3_valid(s2_io_metaReadResp_3_valid),
    .io_metaReadResp_3_dirty(s2_io_metaReadResp_3_dirty),
    .io_dataReadResp_0_data(s2_io_dataReadResp_0_data),
    .io_dataReadResp_1_data(s2_io_dataReadResp_1_data),
    .io_dataReadResp_2_data(s2_io_dataReadResp_2_data),
    .io_dataReadResp_3_data(s2_io_dataReadResp_3_data),
    .io_metaWriteBus_req_valid(s2_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s2_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s2_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_data_dirty(s2_io_metaWriteBus_req_bits_data_dirty),
    .io_metaWriteBus_req_bits_waymask(s2_io_metaWriteBus_req_bits_waymask),
    .io_dataWriteBus_req_valid(s2_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s2_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s2_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s2_io_dataWriteBus_req_bits_waymask),
    .DISPLAY_ENABLE(s2_DISPLAY_ENABLE)
  );
  CacheStage3_2 s3 ( // @[Cache.scala 477:18]
    .clock(s3_clock),
    .reset(s3_reset),
    .io_in_ready(s3_io_in_ready),
    .io_in_valid(s3_io_in_valid),
    .io_in_bits_req_addr(s3_io_in_bits_req_addr),
    .io_in_bits_req_size(s3_io_in_bits_req_size),
    .io_in_bits_req_cmd(s3_io_in_bits_req_cmd),
    .io_in_bits_req_wmask(s3_io_in_bits_req_wmask),
    .io_in_bits_req_wdata(s3_io_in_bits_req_wdata),
    .io_in_bits_metas_0_tag(s3_io_in_bits_metas_0_tag),
    .io_in_bits_metas_0_valid(s3_io_in_bits_metas_0_valid),
    .io_in_bits_metas_0_dirty(s3_io_in_bits_metas_0_dirty),
    .io_in_bits_metas_1_tag(s3_io_in_bits_metas_1_tag),
    .io_in_bits_metas_1_valid(s3_io_in_bits_metas_1_valid),
    .io_in_bits_metas_1_dirty(s3_io_in_bits_metas_1_dirty),
    .io_in_bits_metas_2_tag(s3_io_in_bits_metas_2_tag),
    .io_in_bits_metas_2_valid(s3_io_in_bits_metas_2_valid),
    .io_in_bits_metas_2_dirty(s3_io_in_bits_metas_2_dirty),
    .io_in_bits_metas_3_tag(s3_io_in_bits_metas_3_tag),
    .io_in_bits_metas_3_valid(s3_io_in_bits_metas_3_valid),
    .io_in_bits_metas_3_dirty(s3_io_in_bits_metas_3_dirty),
    .io_in_bits_datas_0_data(s3_io_in_bits_datas_0_data),
    .io_in_bits_datas_1_data(s3_io_in_bits_datas_1_data),
    .io_in_bits_datas_2_data(s3_io_in_bits_datas_2_data),
    .io_in_bits_datas_3_data(s3_io_in_bits_datas_3_data),
    .io_in_bits_hit(s3_io_in_bits_hit),
    .io_in_bits_waymask(s3_io_in_bits_waymask),
    .io_in_bits_mmio(s3_io_in_bits_mmio),
    .io_in_bits_isForwardData(s3_io_in_bits_isForwardData),
    .io_in_bits_forwardData_data_data(s3_io_in_bits_forwardData_data_data),
    .io_in_bits_forwardData_waymask(s3_io_in_bits_forwardData_waymask),
    .io_out_ready(s3_io_out_ready),
    .io_out_valid(s3_io_out_valid),
    .io_out_bits_cmd(s3_io_out_bits_cmd),
    .io_out_bits_rdata(s3_io_out_bits_rdata),
    .io_isFinish(s3_io_isFinish),
    .io_dataReadBus_req_ready(s3_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s3_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s3_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s3_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s3_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s3_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s3_io_dataReadBus_resp_data_3_data),
    .io_dataWriteBus_req_valid(s3_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s3_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s3_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s3_io_dataWriteBus_req_bits_waymask),
    .io_metaWriteBus_req_valid(s3_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s3_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s3_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_data_valid(s3_io_metaWriteBus_req_bits_data_valid),
    .io_metaWriteBus_req_bits_data_dirty(s3_io_metaWriteBus_req_bits_data_dirty),
    .io_metaWriteBus_req_bits_waymask(s3_io_metaWriteBus_req_bits_waymask),
    .io_mem_req_ready(s3_io_mem_req_ready),
    .io_mem_req_valid(s3_io_mem_req_valid),
    .io_mem_req_bits_addr(s3_io_mem_req_bits_addr),
    .io_mem_req_bits_size(s3_io_mem_req_bits_size),
    .io_mem_req_bits_cmd(s3_io_mem_req_bits_cmd),
    .io_mem_req_bits_wmask(s3_io_mem_req_bits_wmask),
    .io_mem_req_bits_wdata(s3_io_mem_req_bits_wdata),
    .io_mem_resp_ready(s3_io_mem_resp_ready),
    .io_mem_resp_valid(s3_io_mem_resp_valid),
    .io_mem_resp_bits_cmd(s3_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_rdata(s3_io_mem_resp_bits_rdata),
    .io_cohResp_valid(s3_io_cohResp_valid),
    .io_dataReadRespToL1(s3_io_dataReadRespToL1),
    .DISPLAY_ENABLE(s3_DISPLAY_ENABLE)
  );
  SRAMTemplateWithArbiter_4 metaArray ( // @[Cache.scala 478:25]
    .clock(metaArray_clock),
    .reset(metaArray_reset),
    .io_r_0_req_ready(metaArray_io_r_0_req_ready),
    .io_r_0_req_valid(metaArray_io_r_0_req_valid),
    .io_r_0_req_bits_setIdx(metaArray_io_r_0_req_bits_setIdx),
    .io_r_0_resp_data_0_tag(metaArray_io_r_0_resp_data_0_tag),
    .io_r_0_resp_data_0_valid(metaArray_io_r_0_resp_data_0_valid),
    .io_r_0_resp_data_0_dirty(metaArray_io_r_0_resp_data_0_dirty),
    .io_r_0_resp_data_1_tag(metaArray_io_r_0_resp_data_1_tag),
    .io_r_0_resp_data_1_valid(metaArray_io_r_0_resp_data_1_valid),
    .io_r_0_resp_data_1_dirty(metaArray_io_r_0_resp_data_1_dirty),
    .io_r_0_resp_data_2_tag(metaArray_io_r_0_resp_data_2_tag),
    .io_r_0_resp_data_2_valid(metaArray_io_r_0_resp_data_2_valid),
    .io_r_0_resp_data_2_dirty(metaArray_io_r_0_resp_data_2_dirty),
    .io_r_0_resp_data_3_tag(metaArray_io_r_0_resp_data_3_tag),
    .io_r_0_resp_data_3_valid(metaArray_io_r_0_resp_data_3_valid),
    .io_r_0_resp_data_3_dirty(metaArray_io_r_0_resp_data_3_dirty),
    .io_w_req_valid(metaArray_io_w_req_valid),
    .io_w_req_bits_setIdx(metaArray_io_w_req_bits_setIdx),
    .io_w_req_bits_data_tag(metaArray_io_w_req_bits_data_tag),
    .io_w_req_bits_data_dirty(metaArray_io_w_req_bits_data_dirty),
    .io_w_req_bits_waymask(metaArray_io_w_req_bits_waymask)
  );
  SRAMTemplateWithArbiter_5 dataArray ( // @[Cache.scala 479:25]
    .clock(dataArray_clock),
    .reset(dataArray_reset),
    .io_r_0_req_ready(dataArray_io_r_0_req_ready),
    .io_r_0_req_valid(dataArray_io_r_0_req_valid),
    .io_r_0_req_bits_setIdx(dataArray_io_r_0_req_bits_setIdx),
    .io_r_0_resp_data_0_data(dataArray_io_r_0_resp_data_0_data),
    .io_r_0_resp_data_1_data(dataArray_io_r_0_resp_data_1_data),
    .io_r_0_resp_data_2_data(dataArray_io_r_0_resp_data_2_data),
    .io_r_0_resp_data_3_data(dataArray_io_r_0_resp_data_3_data),
    .io_r_1_req_ready(dataArray_io_r_1_req_ready),
    .io_r_1_req_valid(dataArray_io_r_1_req_valid),
    .io_r_1_req_bits_setIdx(dataArray_io_r_1_req_bits_setIdx),
    .io_r_1_resp_data_0_data(dataArray_io_r_1_resp_data_0_data),
    .io_r_1_resp_data_1_data(dataArray_io_r_1_resp_data_1_data),
    .io_r_1_resp_data_2_data(dataArray_io_r_1_resp_data_2_data),
    .io_r_1_resp_data_3_data(dataArray_io_r_1_resp_data_3_data),
    .io_w_req_valid(dataArray_io_w_req_valid),
    .io_w_req_bits_setIdx(dataArray_io_w_req_bits_setIdx),
    .io_w_req_bits_data_data(dataArray_io_w_req_bits_data_data),
    .io_w_req_bits_waymask(dataArray_io_w_req_bits_waymask)
  );
  Arbiter_9 arb ( // @[Cache.scala 488:19]
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_addr(arb_io_in_0_bits_addr),
    .io_in_0_bits_size(arb_io_in_0_bits_size),
    .io_in_0_bits_cmd(arb_io_in_0_bits_cmd),
    .io_in_0_bits_wmask(arb_io_in_0_bits_wmask),
    .io_in_0_bits_wdata(arb_io_in_0_bits_wdata),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_addr(arb_io_in_1_bits_addr),
    .io_in_1_bits_size(arb_io_in_1_bits_size),
    .io_in_1_bits_cmd(arb_io_in_1_bits_cmd),
    .io_in_1_bits_wmask(arb_io_in_1_bits_wmask),
    .io_in_1_bits_wdata(arb_io_in_1_bits_wdata),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_addr(arb_io_out_bits_addr),
    .io_out_bits_size(arb_io_out_bits_size),
    .io_out_bits_cmd(arb_io_out_bits_cmd),
    .io_out_bits_wmask(arb_io_out_bits_wmask),
    .io_out_bits_wdata(arb_io_out_bits_wdata)
  );
  assign io_in_req_ready = arb_io_in_1_ready; // @[Cache.scala 489:28]
  assign io_in_resp_valid = _T_16 ? 1'h0 : _T_17; // @[Cache.scala 499:14 Cache.scala 505:20]
  assign io_in_resp_bits_cmd = s3_io_out_bits_cmd; // @[Cache.scala 499:14]
  assign io_in_resp_bits_rdata = s3_io_out_bits_rdata; // @[Cache.scala 499:14]
  assign io_out_mem_req_valid = s3_io_mem_req_valid; // @[Cache.scala 501:14]
  assign io_out_mem_req_bits_addr = s3_io_mem_req_bits_addr; // @[Cache.scala 501:14]
  assign io_out_mem_req_bits_cmd = s3_io_mem_req_bits_cmd; // @[Cache.scala 501:14]
  assign io_out_mem_req_bits_wdata = s3_io_mem_req_bits_wdata; // @[Cache.scala 501:14]
  assign s1_clock = clock;
  assign s1_reset = reset;
  assign s1_io_in_valid = arb_io_out_valid; // @[Cache.scala 491:12]
  assign s1_io_in_bits_addr = arb_io_out_bits_addr; // @[Cache.scala 491:12]
  assign s1_io_in_bits_size = arb_io_out_bits_size; // @[Cache.scala 491:12]
  assign s1_io_in_bits_cmd = arb_io_out_bits_cmd; // @[Cache.scala 491:12]
  assign s1_io_in_bits_wmask = arb_io_out_bits_wmask; // @[Cache.scala 491:12]
  assign s1_io_in_bits_wdata = arb_io_out_bits_wdata; // @[Cache.scala 491:12]
  assign s1_io_out_ready = s2_io_in_ready; // @[Pipeline.scala 29:16]
  assign s1_io_metaReadBus_req_ready = metaArray_io_r_0_req_ready; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_0_tag = metaArray_io_r_0_resp_data_0_tag; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_0_valid = metaArray_io_r_0_resp_data_0_valid; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_0_dirty = metaArray_io_r_0_resp_data_0_dirty; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_1_tag = metaArray_io_r_0_resp_data_1_tag; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_1_valid = metaArray_io_r_0_resp_data_1_valid; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_1_dirty = metaArray_io_r_0_resp_data_1_dirty; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_2_tag = metaArray_io_r_0_resp_data_2_tag; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_2_valid = metaArray_io_r_0_resp_data_2_valid; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_2_dirty = metaArray_io_r_0_resp_data_2_dirty; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_3_tag = metaArray_io_r_0_resp_data_3_tag; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_3_valid = metaArray_io_r_0_resp_data_3_valid; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_3_dirty = metaArray_io_r_0_resp_data_3_dirty; // @[Cache.scala 523:21]
  assign s1_io_dataReadBus_req_ready = dataArray_io_r_0_req_ready; // @[Cache.scala 524:21]
  assign s1_io_dataReadBus_resp_data_0_data = dataArray_io_r_0_resp_data_0_data; // @[Cache.scala 524:21]
  assign s1_io_dataReadBus_resp_data_1_data = dataArray_io_r_0_resp_data_1_data; // @[Cache.scala 524:21]
  assign s1_io_dataReadBus_resp_data_2_data = dataArray_io_r_0_resp_data_2_data; // @[Cache.scala 524:21]
  assign s1_io_dataReadBus_resp_data_3_data = dataArray_io_r_0_resp_data_3_data; // @[Cache.scala 524:21]
  assign s1_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign s2_clock = clock;
  assign s2_reset = reset;
  assign s2_io_in_valid = _T_2; // @[Pipeline.scala 31:17]
  assign s2_io_in_bits_req_addr = _T_5_req_addr; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_size = _T_5_req_size; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_cmd = _T_5_req_cmd; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_wmask = _T_5_req_wmask; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_wdata = _T_5_req_wdata; // @[Pipeline.scala 30:16]
  assign s2_io_out_ready = s3_io_in_ready; // @[Pipeline.scala 29:16]
  assign s2_io_metaReadResp_0_tag = s1_io_metaReadBus_resp_data_0_tag; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_0_valid = s1_io_metaReadBus_resp_data_0_valid; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_0_dirty = s1_io_metaReadBus_resp_data_0_dirty; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_1_tag = s1_io_metaReadBus_resp_data_1_tag; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_1_valid = s1_io_metaReadBus_resp_data_1_valid; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_1_dirty = s1_io_metaReadBus_resp_data_1_dirty; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_2_tag = s1_io_metaReadBus_resp_data_2_tag; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_2_valid = s1_io_metaReadBus_resp_data_2_valid; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_2_dirty = s1_io_metaReadBus_resp_data_2_dirty; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_3_tag = s1_io_metaReadBus_resp_data_3_tag; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_3_valid = s1_io_metaReadBus_resp_data_3_valid; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_3_dirty = s1_io_metaReadBus_resp_data_3_dirty; // @[Cache.scala 530:22]
  assign s2_io_dataReadResp_0_data = s1_io_dataReadBus_resp_data_0_data; // @[Cache.scala 531:22]
  assign s2_io_dataReadResp_1_data = s1_io_dataReadBus_resp_data_1_data; // @[Cache.scala 531:22]
  assign s2_io_dataReadResp_2_data = s1_io_dataReadBus_resp_data_2_data; // @[Cache.scala 531:22]
  assign s2_io_dataReadResp_3_data = s1_io_dataReadBus_resp_data_3_data; // @[Cache.scala 531:22]
  assign s2_io_metaWriteBus_req_valid = s3_io_metaWriteBus_req_valid; // @[Cache.scala 533:22]
  assign s2_io_metaWriteBus_req_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 533:22]
  assign s2_io_metaWriteBus_req_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 533:22]
  assign s2_io_metaWriteBus_req_bits_data_dirty = s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 533:22]
  assign s2_io_metaWriteBus_req_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 533:22]
  assign s2_io_dataWriteBus_req_valid = s3_io_dataWriteBus_req_valid; // @[Cache.scala 532:22]
  assign s2_io_dataWriteBus_req_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 532:22]
  assign s2_io_dataWriteBus_req_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 532:22]
  assign s2_io_dataWriteBus_req_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 532:22]
  assign s2_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign s3_clock = clock;
  assign s3_reset = reset;
  assign s3_io_in_valid = _T_7; // @[Pipeline.scala 31:17]
  assign s3_io_in_bits_req_addr = _T_10_req_addr; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_size = _T_10_req_size; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_cmd = _T_10_req_cmd; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_wmask = _T_10_req_wmask; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_wdata = _T_10_req_wdata; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_tag = _T_10_metas_0_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_valid = _T_10_metas_0_valid; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_dirty = _T_10_metas_0_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_tag = _T_10_metas_1_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_valid = _T_10_metas_1_valid; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_dirty = _T_10_metas_1_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_tag = _T_10_metas_2_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_valid = _T_10_metas_2_valid; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_dirty = _T_10_metas_2_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_tag = _T_10_metas_3_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_valid = _T_10_metas_3_valid; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_dirty = _T_10_metas_3_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_0_data = _T_10_datas_0_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_1_data = _T_10_datas_1_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_2_data = _T_10_datas_2_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_3_data = _T_10_datas_3_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_hit = _T_10_hit; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_waymask = _T_10_waymask; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_mmio = _T_10_mmio; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_isForwardData = _T_10_isForwardData; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_data_data = _T_10_forwardData_data_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_waymask = _T_10_forwardData_waymask; // @[Pipeline.scala 30:16]
  assign s3_io_out_ready = 1'h1; // @[Cache.scala 499:14]
  assign s3_io_dataReadBus_req_ready = dataArray_io_r_1_req_ready; // @[Cache.scala 525:21]
  assign s3_io_dataReadBus_resp_data_0_data = dataArray_io_r_1_resp_data_0_data; // @[Cache.scala 525:21]
  assign s3_io_dataReadBus_resp_data_1_data = dataArray_io_r_1_resp_data_1_data; // @[Cache.scala 525:21]
  assign s3_io_dataReadBus_resp_data_2_data = dataArray_io_r_1_resp_data_2_data; // @[Cache.scala 525:21]
  assign s3_io_dataReadBus_resp_data_3_data = dataArray_io_r_1_resp_data_3_data; // @[Cache.scala 525:21]
  assign s3_io_mem_req_ready = io_out_mem_req_ready; // @[Cache.scala 501:14]
  assign s3_io_mem_resp_valid = io_out_mem_resp_valid; // @[Cache.scala 501:14]
  assign s3_io_mem_resp_bits_cmd = io_out_mem_resp_bits_cmd; // @[Cache.scala 501:14]
  assign s3_io_mem_resp_bits_rdata = io_out_mem_resp_bits_rdata; // @[Cache.scala 501:14]
  assign s3_DISPLAY_ENABLE = DISPLAY_ENABLE;
  assign metaArray_clock = clock;
  assign metaArray_reset = reset;
  assign metaArray_io_r_0_req_valid = s1_io_metaReadBus_req_valid; // @[Cache.scala 523:21]
  assign metaArray_io_r_0_req_bits_setIdx = s1_io_metaReadBus_req_bits_setIdx; // @[Cache.scala 523:21]
  assign metaArray_io_w_req_valid = s3_io_metaWriteBus_req_valid; // @[Cache.scala 527:18]
  assign metaArray_io_w_req_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 527:18]
  assign metaArray_io_w_req_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 527:18]
  assign metaArray_io_w_req_bits_data_dirty = s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 527:18]
  assign metaArray_io_w_req_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 527:18]
  assign dataArray_clock = clock;
  assign dataArray_reset = reset;
  assign dataArray_io_r_0_req_valid = s1_io_dataReadBus_req_valid; // @[Cache.scala 524:21]
  assign dataArray_io_r_0_req_bits_setIdx = s1_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 524:21]
  assign dataArray_io_r_1_req_valid = s3_io_dataReadBus_req_valid; // @[Cache.scala 525:21]
  assign dataArray_io_r_1_req_bits_setIdx = s3_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 525:21]
  assign dataArray_io_w_req_valid = s3_io_dataWriteBus_req_valid; // @[Cache.scala 528:18]
  assign dataArray_io_w_req_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 528:18]
  assign dataArray_io_w_req_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 528:18]
  assign dataArray_io_w_req_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 528:18]
  assign arb_io_in_0_valid = 1'h0; // @[Cache.scala 513:24]
  assign arb_io_in_0_bits_addr = 32'h0; // @[Cache.scala 512:23]
  assign arb_io_in_0_bits_size = 3'h0; // @[Cache.scala 512:23]
  assign arb_io_in_0_bits_cmd = 4'h0; // @[Cache.scala 512:23]
  assign arb_io_in_0_bits_wmask = 8'h0; // @[Cache.scala 512:23]
  assign arb_io_in_0_bits_wdata = 64'h0; // @[Cache.scala 512:23]
  assign arb_io_in_1_valid = io_in_req_valid; // @[Cache.scala 489:28]
  assign arb_io_in_1_bits_addr = io_in_req_bits_addr; // @[Cache.scala 489:28]
  assign arb_io_in_1_bits_size = io_in_req_bits_size; // @[Cache.scala 489:28]
  assign arb_io_in_1_bits_cmd = io_in_req_bits_cmd; // @[Cache.scala 489:28]
  assign arb_io_in_1_bits_wmask = io_in_req_bits_wmask; // @[Cache.scala 489:28]
  assign arb_io_in_1_bits_wdata = io_in_req_bits_wdata; // @[Cache.scala 489:28]
  assign arb_io_out_ready = s1_io_in_ready; // @[Cache.scala 491:12]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _T_5_req_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_5_req_size = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  _T_5_req_cmd = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  _T_5_req_wmask = _RAND_4[7:0];
  _RAND_5 = {2{`RANDOM}};
  _T_5_req_wdata = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  _T_7 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_10_req_addr = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  _T_10_req_size = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  _T_10_req_cmd = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  _T_10_req_wmask = _RAND_10[7:0];
  _RAND_11 = {2{`RANDOM}};
  _T_10_req_wdata = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  _T_10_metas_0_tag = _RAND_12[16:0];
  _RAND_13 = {1{`RANDOM}};
  _T_10_metas_0_valid = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  _T_10_metas_0_dirty = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  _T_10_metas_1_tag = _RAND_15[16:0];
  _RAND_16 = {1{`RANDOM}};
  _T_10_metas_1_valid = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  _T_10_metas_1_dirty = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  _T_10_metas_2_tag = _RAND_18[16:0];
  _RAND_19 = {1{`RANDOM}};
  _T_10_metas_2_valid = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  _T_10_metas_2_dirty = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  _T_10_metas_3_tag = _RAND_21[16:0];
  _RAND_22 = {1{`RANDOM}};
  _T_10_metas_3_valid = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  _T_10_metas_3_dirty = _RAND_23[0:0];
  _RAND_24 = {2{`RANDOM}};
  _T_10_datas_0_data = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  _T_10_datas_1_data = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  _T_10_datas_2_data = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  _T_10_datas_3_data = _RAND_27[63:0];
  _RAND_28 = {1{`RANDOM}};
  _T_10_hit = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  _T_10_waymask = _RAND_29[3:0];
  _RAND_30 = {1{`RANDOM}};
  _T_10_mmio = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  _T_10_isForwardData = _RAND_31[0:0];
  _RAND_32 = {2{`RANDOM}};
  _T_10_forwardData_data_data = _RAND_32[63:0];
  _RAND_33 = {1{`RANDOM}};
  _T_10_forwardData_waymask = _RAND_33[3:0];
  _RAND_34 = {2{`RANDOM}};
  _T_20 = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  _T_29 = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  _T_38 = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  _T_47 = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  _T_56 = _RAND_38[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_2 <= 1'h0;
    end else begin
      _T_2 <= _GEN_1;
    end
    if (_T_3) begin
      _T_5_req_addr <= s1_io_out_bits_req_addr;
    end
    if (_T_3) begin
      _T_5_req_size <= s1_io_out_bits_req_size;
    end
    if (_T_3) begin
      _T_5_req_cmd <= s1_io_out_bits_req_cmd;
    end
    if (_T_3) begin
      _T_5_req_wmask <= s1_io_out_bits_req_wmask;
    end
    if (_T_3) begin
      _T_5_req_wdata <= s1_io_out_bits_req_wdata;
    end
    if (reset) begin
      _T_7 <= 1'h0;
    end else begin
      _T_7 <= _GEN_9;
    end
    if (_T_8) begin
      _T_10_req_addr <= s2_io_out_bits_req_addr;
    end
    if (_T_8) begin
      _T_10_req_size <= s2_io_out_bits_req_size;
    end
    if (_T_8) begin
      _T_10_req_cmd <= s2_io_out_bits_req_cmd;
    end
    if (_T_8) begin
      _T_10_req_wmask <= s2_io_out_bits_req_wmask;
    end
    if (_T_8) begin
      _T_10_req_wdata <= s2_io_out_bits_req_wdata;
    end
    if (_T_8) begin
      _T_10_metas_0_tag <= s2_io_out_bits_metas_0_tag;
    end
    if (_T_8) begin
      _T_10_metas_0_valid <= s2_io_out_bits_metas_0_valid;
    end
    if (_T_8) begin
      _T_10_metas_0_dirty <= s2_io_out_bits_metas_0_dirty;
    end
    if (_T_8) begin
      _T_10_metas_1_tag <= s2_io_out_bits_metas_1_tag;
    end
    if (_T_8) begin
      _T_10_metas_1_valid <= s2_io_out_bits_metas_1_valid;
    end
    if (_T_8) begin
      _T_10_metas_1_dirty <= s2_io_out_bits_metas_1_dirty;
    end
    if (_T_8) begin
      _T_10_metas_2_tag <= s2_io_out_bits_metas_2_tag;
    end
    if (_T_8) begin
      _T_10_metas_2_valid <= s2_io_out_bits_metas_2_valid;
    end
    if (_T_8) begin
      _T_10_metas_2_dirty <= s2_io_out_bits_metas_2_dirty;
    end
    if (_T_8) begin
      _T_10_metas_3_tag <= s2_io_out_bits_metas_3_tag;
    end
    if (_T_8) begin
      _T_10_metas_3_valid <= s2_io_out_bits_metas_3_valid;
    end
    if (_T_8) begin
      _T_10_metas_3_dirty <= s2_io_out_bits_metas_3_dirty;
    end
    if (_T_8) begin
      _T_10_datas_0_data <= s2_io_out_bits_datas_0_data;
    end
    if (_T_8) begin
      _T_10_datas_1_data <= s2_io_out_bits_datas_1_data;
    end
    if (_T_8) begin
      _T_10_datas_2_data <= s2_io_out_bits_datas_2_data;
    end
    if (_T_8) begin
      _T_10_datas_3_data <= s2_io_out_bits_datas_3_data;
    end
    if (_T_8) begin
      _T_10_hit <= s2_io_out_bits_hit;
    end
    if (_T_8) begin
      _T_10_waymask <= s2_io_out_bits_waymask;
    end
    if (_T_8) begin
      _T_10_mmio <= s2_io_out_bits_mmio;
    end
    if (_T_8) begin
      _T_10_isForwardData <= s2_io_out_bits_isForwardData;
    end
    if (_T_8) begin
      _T_10_forwardData_data_data <= s2_io_out_bits_forwardData_data_data;
    end
    if (_T_8) begin
      _T_10_forwardData_waymask <= s2_io_out_bits_forwardData_waymask;
    end
    if (reset) begin
      _T_20 <= 64'h0;
    end else begin
      _T_20 <= _T_22;
    end
    if (reset) begin
      _T_29 <= 64'h0;
    end else begin
      _T_29 <= _T_31;
    end
    if (reset) begin
      _T_38 <= 64'h0;
    end else begin
      _T_38 <= _T_40;
    end
    if (reset) begin
      _T_47 <= 64'h0;
    end else begin
      _T_47 <= _T_49;
    end
    if (reset) begin
      _T_56 <= 64'h0;
    end else begin
      _T_56 <= _T_58;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_26) begin
          $fwrite(32'h80000002,"[%d] Cache_2: ",_T_20); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_26) begin
          $fwrite(32'h80000002,"InReq(%d, %d) InResp(%d, %d) \n",io_in_req_valid,io_in_req_ready,io_in_resp_valid,1'h1); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_26) begin
          $fwrite(32'h80000002,"[%d] Cache_2: ",_T_29); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (DISPLAY_ENABLE & _T_26) begin
          $fwrite(32'h80000002,"{IN s1:(%d,%d), s2:(%d,%d), s3:(%d,%d)} {OUT s1:(%d,%d), s2:(%d,%d), s3:(%d,%d)}\n",s1_io_in_valid,s1_io_in_ready,s2_io_in_valid,s2_io_in_ready,s3_io_in_valid,s3_io_in_ready,s1_io_out_valid,s1_io_out_ready,s2_io_out_valid,s2_io_out_ready,s3_io_out_valid,s3_io_out_ready); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_39 & _T_26) begin
          $fwrite(32'h80000002,"[%d] Cache_2: ",_T_38); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_39 & _T_26) begin
          $fwrite(32'h80000002,"[l2cache.S1]: addr = 0x%x, cmd = %d, size = %d, wmask = 0x%x, wdata = 0x%x\n",s1_io_in_bits_addr,s1_io_in_bits_cmd,s1_io_in_bits_size,s1_io_in_bits_wmask,s1_io_in_bits_wdata); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_26) begin
          $fwrite(32'h80000002,"[%d] Cache_2: ",_T_47); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_26) begin
          $fwrite(32'h80000002,"[l2cache.S2]: addr = 0x%x, cmd = %d, size = %d, wmask = 0x%x, wdata = 0x%x\n",s2_io_in_bits_req_addr,s2_io_in_bits_req_cmd,s2_io_in_bits_req_size,s2_io_in_bits_req_wmask,s2_io_in_bits_req_wdata); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_43 & _T_26) begin
          $fwrite(32'h80000002,"[%d] Cache_2: ",_T_56); // @[Debug.scala 56:24]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_43 & _T_26) begin
          $fwrite(32'h80000002,"[l2cache.S3]: addr = 0x%x, cmd = %d, size = %d, wmask = 0x%x, wdata = 0x%x\n",s3_io_in_bits_req_addr,s3_io_in_bits_req_cmd,s3_io_in_bits_req_size,s3_io_in_bits_req_wmask,s3_io_in_bits_req_wdata); // @[Debug.scala 57:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module SimpleBusAddressMapper(
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [3:0]  io_in_req_bits_cmd,
  input  [63:0] io_in_req_bits_wdata,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [3:0]  io_out_req_bits_cmd,
  output [63:0] io_out_req_bits_wdata,
  input         io_out_resp_valid,
  input  [3:0]  io_out_resp_bits_cmd,
  input  [63:0] io_out_resp_bits_rdata
);
  assign io_in_req_ready = io_out_req_ready; // @[AddressMapper.scala 31:10]
  assign io_in_resp_valid = io_out_resp_valid; // @[AddressMapper.scala 31:10]
  assign io_in_resp_bits_cmd = io_out_resp_bits_cmd; // @[AddressMapper.scala 31:10]
  assign io_in_resp_bits_rdata = io_out_resp_bits_rdata; // @[AddressMapper.scala 31:10]
  assign io_out_req_valid = io_in_req_valid; // @[AddressMapper.scala 31:10]
  assign io_out_req_bits_addr = io_in_req_bits_addr; // @[AddressMapper.scala 31:10]
  assign io_out_req_bits_cmd = io_in_req_bits_cmd; // @[AddressMapper.scala 31:10]
  assign io_out_req_bits_wdata = io_in_req_bits_wdata; // @[AddressMapper.scala 31:10]
endmodule
module SimpleBus2AXI4Converter(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [3:0]  io_in_req_bits_cmd,
  input  [63:0] io_in_req_bits_wdata,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_aw_ready,
  output        io_out_aw_valid,
  output [31:0] io_out_aw_bits_addr,
  output [7:0]  io_out_aw_bits_len,
  output [2:0]  io_out_aw_bits_size,
  output [1:0]  io_out_aw_bits_burst,
  input         io_out_w_ready,
  output        io_out_w_valid,
  output [63:0] io_out_w_bits_data,
  output        io_out_w_bits_last,
  input         io_out_b_valid,
  input         io_out_ar_ready,
  output        io_out_ar_valid,
  output [31:0] io_out_ar_bits_addr,
  output [7:0]  io_out_ar_bits_len,
  output [2:0]  io_out_ar_bits_size,
  output [1:0]  io_out_ar_bits_burst,
  input         io_out_r_valid,
  input  [63:0] io_out_r_bits_data,
  input         io_out_r_bits_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] _T_8 = io_in_req_bits_cmd[1] ? 3'h7 : 3'h0; // @[ToAXI4.scala 169:30]
  wire  _T_9 = io_in_req_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_10 = io_in_req_bits_cmd == 4'h1; // @[SimpleBus.scala 77:29]
  wire [2:0] _T_12 = io_out_r_bits_last ? 3'h6 : 3'h0; // @[ToAXI4.scala 184:28]
  wire  _T_13 = io_out_aw_ready & io_out_aw_valid; // @[Decoupled.scala 40:37]
  reg  awAck; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_13 | awAck; // @[StopWatch.scala 30:20]
  wire  _T_17 = io_out_w_ready & io_out_w_valid; // @[Decoupled.scala 40:37]
  wire  _T_18 = _T_13 & _T_17; // @[ToAXI4.scala 189:27]
  wire  _T_19 = _T_18 & io_out_w_bits_last; // @[ToAXI4.scala 189:43]
  reg  wAck; // @[StopWatch.scala 24:20]
  wire  _T_20 = awAck & wAck; // @[ToAXI4.scala 189:63]
  wire  wSend = _T_19 | _T_20; // @[ToAXI4.scala 189:53]
  wire  _T_15 = _T_17 & io_out_w_bits_last; // @[ToAXI4.scala 188:41]
  wire  _GEN_2 = _T_15 | wAck; // @[StopWatch.scala 30:20]
  wire  _T_23 = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 40:37]
  reg  wen; // @[Reg.scala 15:16]
  wire  _T_25 = ~io_in_req_bits_cmd[0]; // @[SimpleBus.scala 73:18]
  wire  _T_27 = ~io_in_req_bits_cmd[3]; // @[SimpleBus.scala 73:29]
  wire  _T_28 = _T_25 & _T_27; // @[SimpleBus.scala 73:26]
  wire  _T_31 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[SimpleBus.scala 103:29]
  wire  _T_32 = ~awAck; // @[ToAXI4.scala 193:36]
  wire  _T_36 = ~wAck; // @[ToAXI4.scala 194:36]
  wire  _T_40 = _T_36 & io_out_w_ready; // @[ToAXI4.scala 195:55]
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _T_40 : io_out_ar_ready; // @[ToAXI4.scala 195:18]
  assign io_in_resp_valid = wen ? io_out_b_valid : io_out_r_valid; // @[ToAXI4.scala 199:19]
  assign io_in_resp_bits_cmd = {{1'd0}, _T_12}; // @[ToAXI4.scala 184:22]
  assign io_in_resp_bits_rdata = io_out_r_bits_data; // @[ToAXI4.scala 183:23]
  assign io_out_aw_valid = _T_31 & _T_32; // @[ToAXI4.scala 193:16]
  assign io_out_aw_bits_addr = io_out_ar_bits_addr; // @[ToAXI4.scala 182:6]
  assign io_out_aw_bits_len = io_out_ar_bits_len; // @[ToAXI4.scala 182:6]
  assign io_out_aw_bits_size = io_out_ar_bits_size; // @[ToAXI4.scala 182:6]
  assign io_out_aw_bits_burst = io_out_ar_bits_burst; // @[ToAXI4.scala 182:6]
  assign io_out_w_valid = _T_31 & _T_36; // @[ToAXI4.scala 194:16]
  assign io_out_w_bits_data = io_in_req_bits_wdata; // @[ToAXI4.scala 160:10]
  assign io_out_w_bits_last = _T_9 | _T_10; // @[ToAXI4.scala 177:24]
  assign io_out_ar_valid = io_in_req_valid & _T_28; // @[ToAXI4.scala 192:16]
  assign io_out_ar_bits_addr = io_in_req_bits_addr; // @[ToAXI4.scala 158:12]
  assign io_out_ar_bits_len = {{5'd0}, _T_8}; // @[ToAXI4.scala 169:24]
  assign io_out_ar_bits_size = 3'h3; // @[ToAXI4.scala 170:24]
  assign io_out_ar_bits_burst = 2'h2; // @[ToAXI4.scala 171:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  awAck = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wAck = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wen = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      awAck <= 1'h0;
    end else if (wSend) begin
      awAck <= 1'h0;
    end else begin
      awAck <= _GEN_0;
    end
    if (reset) begin
      wAck <= 1'h0;
    end else if (wSend) begin
      wAck <= 1'h0;
    end else begin
      wAck <= _GEN_2;
    end
    if (_T_23) begin
      wen <= io_in_req_bits_cmd[0];
    end
  end
endmodule
module SimpleBusCrossbar1toN(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [2:0]  io_in_req_bits_size,
  input  [3:0]  io_in_req_bits_cmd,
  input  [7:0]  io_in_req_bits_wmask,
  input  [63:0] io_in_req_bits_wdata,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_0_req_ready,
  output        io_out_0_req_valid,
  output [31:0] io_out_0_req_bits_addr,
  output [2:0]  io_out_0_req_bits_size,
  output [3:0]  io_out_0_req_bits_cmd,
  output [7:0]  io_out_0_req_bits_wmask,
  output [63:0] io_out_0_req_bits_wdata,
  output        io_out_0_resp_ready,
  input         io_out_0_resp_valid,
  input  [63:0] io_out_0_resp_bits_rdata,
  input         io_out_1_req_ready,
  output        io_out_1_req_valid,
  output [31:0] io_out_1_req_bits_addr,
  output [2:0]  io_out_1_req_bits_size,
  output [3:0]  io_out_1_req_bits_cmd,
  output [7:0]  io_out_1_req_bits_wmask,
  output [63:0] io_out_1_req_bits_wdata,
  output        io_out_1_resp_ready,
  input         io_out_1_resp_valid,
  input  [63:0] io_out_1_resp_bits_rdata,
  input         io_out_2_req_ready,
  output        io_out_2_req_valid,
  output [31:0] io_out_2_req_bits_addr,
  output [2:0]  io_out_2_req_bits_size,
  output [3:0]  io_out_2_req_bits_cmd,
  output [7:0]  io_out_2_req_bits_wmask,
  output [63:0] io_out_2_req_bits_wdata,
  output        io_out_2_resp_ready,
  input         io_out_2_resp_valid,
  input  [63:0] io_out_2_resp_bits_rdata,
  input         DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[Crossbar.scala 31:22]
  wire  _T = io_in_req_bits_addr >= 32'h40000000; // @[Crossbar.scala 36:20]
  wire  _T_1 = io_in_req_bits_addr < 32'h80000000; // @[Crossbar.scala 36:42]
  wire  outSelVec_0 = _T & _T_1; // @[Crossbar.scala 36:34]
  wire  _T_3 = io_in_req_bits_addr >= 32'h38000000; // @[Crossbar.scala 36:20]
  wire  _T_4 = io_in_req_bits_addr < 32'h38010000; // @[Crossbar.scala 36:42]
  wire  outSelVec_1 = _T_3 & _T_4; // @[Crossbar.scala 36:34]
  wire  _T_6 = io_in_req_bits_addr >= 32'h3c000000; // @[Crossbar.scala 36:20]
  wire  _T_7 = io_in_req_bits_addr < 32'h40000000; // @[Crossbar.scala 36:42]
  wire  outSelVec_2 = _T_6 & _T_7; // @[Crossbar.scala 36:34]
  wire [1:0] _T_9 = outSelVec_1 ? 2'h1 : 2'h2; // @[Mux.scala 47:69]
  wire [1:0] outSelIdx = outSelVec_0 ? 2'h0 : _T_9; // @[Mux.scala 47:69]
  wire  _GEN_11 = 2'h1 == outSelIdx ? io_out_1_req_ready : io_out_0_req_ready; // @[Decoupled.scala 40:37]
  wire  _GEN_12 = 2'h1 == outSelIdx ? io_out_1_req_valid : io_out_0_req_valid; // @[Decoupled.scala 40:37]
  wire [31:0] _GEN_13 = 2'h1 == outSelIdx ? io_out_1_req_bits_addr : io_out_0_req_bits_addr; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_14 = 2'h1 == outSelIdx ? io_out_1_req_bits_size : io_out_0_req_bits_size; // @[Decoupled.scala 40:37]
  wire [3:0] _GEN_15 = 2'h1 == outSelIdx ? io_out_1_req_bits_cmd : io_out_0_req_bits_cmd; // @[Decoupled.scala 40:37]
  wire [7:0] _GEN_16 = 2'h1 == outSelIdx ? io_out_1_req_bits_wmask : io_out_0_req_bits_wmask; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_17 = 2'h1 == outSelIdx ? io_out_1_req_bits_wdata : io_out_0_req_bits_wdata; // @[Decoupled.scala 40:37]
  wire  _GEN_18 = 2'h1 == outSelIdx ? io_out_1_resp_ready : io_out_0_resp_ready; // @[Decoupled.scala 40:37]
  wire  _GEN_19 = 2'h1 == outSelIdx ? io_out_1_resp_valid : io_out_0_resp_valid; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_21 = 2'h1 == outSelIdx ? io_out_1_resp_bits_rdata : io_out_0_resp_bits_rdata; // @[Decoupled.scala 40:37]
  wire  _GEN_22 = 2'h2 == outSelIdx ? io_out_2_req_ready : _GEN_11; // @[Decoupled.scala 40:37]
  wire  _GEN_23 = 2'h2 == outSelIdx ? io_out_2_req_valid : _GEN_12; // @[Decoupled.scala 40:37]
  wire [31:0] _GEN_24 = 2'h2 == outSelIdx ? io_out_2_req_bits_addr : _GEN_13; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_25 = 2'h2 == outSelIdx ? io_out_2_req_bits_size : _GEN_14; // @[Decoupled.scala 40:37]
  wire [3:0] _GEN_26 = 2'h2 == outSelIdx ? io_out_2_req_bits_cmd : _GEN_15; // @[Decoupled.scala 40:37]
  wire [7:0] _GEN_27 = 2'h2 == outSelIdx ? io_out_2_req_bits_wmask : _GEN_16; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_28 = 2'h2 == outSelIdx ? io_out_2_req_bits_wdata : _GEN_17; // @[Decoupled.scala 40:37]
  wire  _GEN_29 = 2'h2 == outSelIdx ? io_out_2_resp_ready : _GEN_18; // @[Decoupled.scala 40:37]
  wire  _GEN_30 = 2'h2 == outSelIdx ? io_out_2_resp_valid : _GEN_19; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_32 = 2'h2 == outSelIdx ? io_out_2_resp_bits_rdata : _GEN_21; // @[Decoupled.scala 40:37]
  wire  _T_10 = _GEN_22 & _GEN_23; // @[Decoupled.scala 40:37]
  wire  _T_11 = state == 2'h0; // @[Crossbar.scala 39:72]
  wire  _T_12 = _T_10 & _T_11; // @[Crossbar.scala 39:62]
  reg [1:0] outSelIdxResp; // @[Reg.scala 15:16]
  wire [2:0] _T_14 = {outSelVec_2,outSelVec_1,outSelVec_0}; // @[Crossbar.scala 41:54]
  wire  _T_15 = |_T_14; // @[Crossbar.scala 41:61]
  wire  _T_16 = ~_T_15; // @[Crossbar.scala 41:43]
  wire  reqInvalidAddr = io_in_req_valid & _T_16; // @[Crossbar.scala 41:40]
  wire  _T_24 = &_T_14; // @[Crossbar.scala 43:91]
  wire  _T_25 = io_in_req_valid & _T_24; // @[Crossbar.scala 43:71]
  wire  _T_26 = reqInvalidAddr | _T_25; // @[Crossbar.scala 43:51]
  reg [63:0] _T_29; // @[GTimer.scala 24:20]
  wire [63:0] _T_31 = _T_29 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_33 = ~reset; // @[Crossbar.scala 45:13]
  wire  _T_38 = ~_T_25; // @[Crossbar.scala 49:10]
  wire  _T_40 = _T_38 | reset; // @[Crossbar.scala 49:9]
  wire  _T_41 = ~_T_40; // @[Crossbar.scala 49:9]
  wire  _T_43 = io_in_req_valid & _T_11; // @[Crossbar.scala 54:42]
  wire  _T_51 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_53 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _GEN_54 = 2'h1 == outSelIdxResp ? io_out_1_resp_ready : io_out_0_resp_ready; // @[Decoupled.scala 40:37]
  wire  _GEN_55 = 2'h1 == outSelIdxResp ? io_out_1_resp_valid : io_out_0_resp_valid; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_57 = 2'h1 == outSelIdxResp ? io_out_1_resp_bits_rdata : io_out_0_resp_bits_rdata; // @[Decoupled.scala 40:37]
  wire  _GEN_65 = 2'h2 == outSelIdxResp ? io_out_2_resp_ready : _GEN_54; // @[Decoupled.scala 40:37]
  wire  _GEN_66 = 2'h2 == outSelIdxResp ? io_out_2_resp_valid : _GEN_55; // @[Decoupled.scala 40:37]
  wire  _T_54 = _GEN_65 & _GEN_66; // @[Decoupled.scala 40:37]
  wire  _T_55 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_58 = state == 2'h2; // @[Crossbar.scala 67:55]
  wire  _GEN_77 = 2'h0 == outSelIdxResp; // @[Crossbar.scala 70:25]
  wire  _GEN_78 = 2'h1 == outSelIdxResp; // @[Crossbar.scala 70:25]
  wire  _GEN_79 = 2'h2 == outSelIdxResp; // @[Crossbar.scala 70:25]
  wire  _T_64 = _T_11 & io_in_req_valid; // @[Crossbar.scala 74:28]
  reg [63:0] _T_65; // @[GTimer.scala 24:20]
  wire [63:0] _T_67 = _T_65 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_71; // @[GTimer.scala 24:20]
  wire [63:0] _T_73 = _T_71 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_76 = _GEN_29 & _GEN_30; // @[Decoupled.scala 40:37]
  reg [63:0] _T_77; // @[GTimer.scala 24:20]
  wire [63:0] _T_79 = _T_77 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_83; // @[GTimer.scala 24:20]
  wire [63:0] _T_85 = _T_83 + 64'h1; // @[GTimer.scala 25:12]
  wire  _GEN_83 = _T_26 & DISPLAY_ENABLE; // @[Crossbar.scala 45:13]
  wire  _GEN_84 = DISPLAY_ENABLE & _T_64; // @[Crossbar.scala 75:13]
  wire  _GEN_85 = DISPLAY_ENABLE & _T_10; // @[Crossbar.scala 79:13]
  wire  _GEN_86 = DISPLAY_ENABLE & _T_76; // @[Crossbar.scala 82:13]
  wire  _GEN_87 = DISPLAY_ENABLE & io_in_resp_valid; // @[Crossbar.scala 86:13]
  assign io_in_req_ready = _GEN_22 | reqInvalidAddr; // @[Crossbar.scala 71:19]
  assign io_in_resp_valid = _T_54 | _T_58; // @[Crossbar.scala 67:20]
  assign io_in_resp_bits_cmd = 4'h6; // @[Crossbar.scala 68:19]
  assign io_in_resp_bits_rdata = 2'h2 == outSelIdxResp ? io_out_2_resp_bits_rdata : _GEN_57; // @[Crossbar.scala 68:19]
  assign io_out_0_req_valid = outSelVec_0 & _T_43; // @[Crossbar.scala 54:17]
  assign io_out_0_req_bits_addr = io_in_req_bits_addr; // @[Crossbar.scala 53:16]
  assign io_out_0_req_bits_size = io_in_req_bits_size; // @[Crossbar.scala 53:16]
  assign io_out_0_req_bits_cmd = io_in_req_bits_cmd; // @[Crossbar.scala 53:16]
  assign io_out_0_req_bits_wmask = io_in_req_bits_wmask; // @[Crossbar.scala 53:16]
  assign io_out_0_req_bits_wdata = io_in_req_bits_wdata; // @[Crossbar.scala 53:16]
  assign io_out_0_resp_ready = _GEN_77 | outSelVec_0; // @[Crossbar.scala 55:18 Crossbar.scala 70:25]
  assign io_out_1_req_valid = outSelVec_1 & _T_43; // @[Crossbar.scala 54:17]
  assign io_out_1_req_bits_addr = io_in_req_bits_addr; // @[Crossbar.scala 53:16]
  assign io_out_1_req_bits_size = io_in_req_bits_size; // @[Crossbar.scala 53:16]
  assign io_out_1_req_bits_cmd = io_in_req_bits_cmd; // @[Crossbar.scala 53:16]
  assign io_out_1_req_bits_wmask = io_in_req_bits_wmask; // @[Crossbar.scala 53:16]
  assign io_out_1_req_bits_wdata = io_in_req_bits_wdata; // @[Crossbar.scala 53:16]
  assign io_out_1_resp_ready = _GEN_78 | outSelVec_1; // @[Crossbar.scala 55:18 Crossbar.scala 70:25]
  assign io_out_2_req_valid = outSelVec_2 & _T_43; // @[Crossbar.scala 54:17]
  assign io_out_2_req_bits_addr = io_in_req_bits_addr; // @[Crossbar.scala 53:16]
  assign io_out_2_req_bits_size = io_in_req_bits_size; // @[Crossbar.scala 53:16]
  assign io_out_2_req_bits_cmd = io_in_req_bits_cmd; // @[Crossbar.scala 53:16]
  assign io_out_2_req_bits_wmask = io_in_req_bits_wmask; // @[Crossbar.scala 53:16]
  assign io_out_2_req_bits_wdata = io_in_req_bits_wdata; // @[Crossbar.scala 53:16]
  assign io_out_2_resp_ready = _GEN_79 | outSelVec_2; // @[Crossbar.scala 55:18 Crossbar.scala 70:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  outSelIdxResp = _RAND_1[1:0];
  _RAND_2 = {2{`RANDOM}};
  _T_29 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  _T_65 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  _T_71 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  _T_77 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  _T_83 = _RAND_6[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else if (_T_51) begin
      if (reqInvalidAddr) begin
        state <= 2'h2;
      end else if (_T_10) begin
        state <= 2'h1;
      end
    end else if (_T_53) begin
      if (_T_54) begin
        state <= 2'h0;
      end
    end else if (_T_55) begin
      if (io_in_resp_valid) begin
        state <= 2'h0;
      end
    end
    if (_T_12) begin
      if (outSelVec_0) begin
        outSelIdxResp <= 2'h0;
      end else if (outSelVec_1) begin
        outSelIdxResp <= 2'h1;
      end else begin
        outSelIdxResp <= 2'h2;
      end
    end
    if (reset) begin
      _T_29 <= 64'h0;
    end else begin
      _T_29 <= _T_31;
    end
    if (reset) begin
      _T_65 <= 64'h0;
    end else begin
      _T_65 <= _T_67;
    end
    if (reset) begin
      _T_71 <= 64'h0;
    end else begin
      _T_71 <= _T_73;
    end
    if (reset) begin
      _T_77 <= 64'h0;
    end else begin
      _T_77 <= _T_79;
    end
    if (reset) begin
      _T_83 <= 64'h0;
    end else begin
      _T_83 <= _T_85;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_83 & _T_33) begin
          $fwrite(32'h80000002,"crossbar access bad addr %x, time %d\n",io_in_req_bits_addr,_T_29); // @[Crossbar.scala 45:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_41) begin
          $fwrite(32'h80000002,"Assertion failed: address decode error, bad addr = 0x%x\n\n    at Crossbar.scala:49 assert(!(io.in.req.valid && outSelVec.asUInt.andR), \"address decode error, bad addr = 0x%%x\\n\", addr)\n",io_in_req_bits_addr); // @[Crossbar.scala 49:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_41) begin
          $fatal; // @[Crossbar.scala 49:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_84 & _T_33) begin
          $fwrite(32'h80000002,"%d: xbar: in.req: addr = 0x%x, cmd = %d, size = %d, wmask = 0x%x, wdata = 0x%x\n",_T_65,io_in_req_bits_addr,io_in_req_bits_cmd,io_in_req_bits_size,io_in_req_bits_wmask,io_in_req_bits_wdata); // @[Crossbar.scala 75:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_33) begin
          $fwrite(32'h80000002,"%d: xbar: outSelIdx = %d, outSel.req: addr = 0x%x, cmd = %d, size = %d, wmask = 0x%x, wdata = 0x%x\n",_T_71,outSelIdx,_GEN_24,_GEN_26,_GEN_25,_GEN_27,_GEN_28); // @[Crossbar.scala 79:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_86 & _T_33) begin
          $fwrite(32'h80000002,"%d: xbar: outSelIdx= %d, outSel.resp: rdata = %x, cmd = %d\n",_T_77,outSelIdx,_GEN_32,4'h6); // @[Crossbar.scala 82:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_87 & _T_33) begin
          $fwrite(32'h80000002,"%d: xbar: in.resp: rdata = %x, cmd = %d\n",_T_83,io_in_resp_bits_rdata,io_in_resp_bits_cmd); // @[Crossbar.scala 86:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module AXI4CLINT(
  input         clock,
  input         reset,
  output        io__in_aw_ready,
  input         io__in_aw_valid,
  input  [31:0] io__in_aw_bits_addr,
  output        io__in_w_ready,
  input         io__in_w_valid,
  input  [63:0] io__in_w_bits_data,
  input  [7:0]  io__in_w_bits_strb,
  input         io__in_b_ready,
  output        io__in_b_valid,
  output        io__in_ar_ready,
  input         io__in_ar_valid,
  input  [31:0] io__in_ar_bits_addr,
  input         io__in_r_ready,
  output        io__in_r_valid,
  output [63:0] io__in_r_bits_data,
  output        io__extra_mtip,
  output        io__extra_msip,
  output        io_extra_mtip,
  input         isWFI,
  output        io_extra_msip
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] _T_9 = io__in_w_bits_strb[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_11 = io__in_w_bits_strb[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_13 = io__in_w_bits_strb[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_15 = io__in_w_bits_strb[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_17 = io__in_w_bits_strb[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_19 = io__in_w_bits_strb[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_21 = io__in_w_bits_strb[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_23 = io__in_w_bits_strb[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] fullMask = {_T_23,_T_21,_T_19,_T_17,_T_15,_T_13,_T_11,_T_9}; // @[Cat.scala 29:58]
  wire  _T_30 = io__in_ar_ready & io__in_ar_valid; // @[Decoupled.scala 40:37]
  wire  _T_31 = io__in_r_ready & io__in_r_valid; // @[Decoupled.scala 40:37]
  reg  r_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_31 ? 1'h0 : r_busy; // @[StopWatch.scala 26:19]
  wire  _GEN_1 = _T_30 | _GEN_0; // @[StopWatch.scala 27:20]
  wire  _T_33 = ~r_busy; // @[AXI4Slave.scala 71:32]
  reg  ren; // @[AXI4Slave.scala 73:17]
  wire  _T_42 = _T_30 | r_busy; // @[AXI4Slave.scala 74:52]
  wire  _T_43 = ren & _T_42; // @[AXI4Slave.scala 74:35]
  reg  _T_45; // @[StopWatch.scala 24:20]
  wire  _GEN_2 = _T_31 ? 1'h0 : _T_45; // @[StopWatch.scala 26:19]
  wire  _GEN_3 = _T_43 | _GEN_2; // @[StopWatch.scala 27:20]
  wire  _T_46 = io__in_aw_ready & io__in_aw_valid; // @[Decoupled.scala 40:37]
  wire  _T_47 = io__in_b_ready & io__in_b_valid; // @[Decoupled.scala 40:37]
  reg  w_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_4 = _T_47 ? 1'h0 : w_busy; // @[StopWatch.scala 26:19]
  wire  _GEN_5 = _T_46 | _GEN_4; // @[StopWatch.scala 27:20]
  wire  _T_50 = io__in_w_ready & io__in_w_valid; // @[Decoupled.scala 40:37]
  reg  _T_53; // @[StopWatch.scala 24:20]
  wire  _GEN_6 = _T_47 ? 1'h0 : _T_53; // @[StopWatch.scala 26:19]
  wire  _GEN_7 = _T_50 | _GEN_6; // @[StopWatch.scala 27:20]
  reg [63:0] mtime; // @[AXI4CLINT.scala 32:22]
  reg [63:0] mtimecmp; // @[AXI4CLINT.scala 33:25]
  reg [63:0] msip; // @[AXI4CLINT.scala 34:21]
  reg [15:0] freq; // @[AXI4CLINT.scala 37:21]
  reg [15:0] inc; // @[AXI4CLINT.scala 38:20]
  reg [15:0] cnt; // @[AXI4CLINT.scala 40:20]
  wire [15:0] nextCnt = cnt + 16'h1; // @[AXI4CLINT.scala 41:21]
  wire  _T_55 = nextCnt < freq; // @[AXI4CLINT.scala 42:22]
  wire  tick = nextCnt == freq; // @[AXI4CLINT.scala 43:23]
  wire [63:0] _GEN_15 = {{48'd0}, inc}; // @[AXI4CLINT.scala 44:32]
  wire [63:0] _T_58 = mtime + _GEN_15; // @[AXI4CLINT.scala 44:32]
  wire [63:0] _T_61 = mtime + 64'h186a0; // @[AXI4CLINT.scala 49:35]
  wire  _T_96 = 16'h0 == io__in_ar_bits_addr[15:0]; // @[LookupTree.scala 24:34]
  wire  _T_97 = 16'h8000 == io__in_ar_bits_addr[15:0]; // @[LookupTree.scala 24:34]
  wire  _T_98 = 16'hbff8 == io__in_ar_bits_addr[15:0]; // @[LookupTree.scala 24:34]
  wire  _T_99 = 16'h8008 == io__in_ar_bits_addr[15:0]; // @[LookupTree.scala 24:34]
  wire  _T_100 = 16'h4000 == io__in_ar_bits_addr[15:0]; // @[LookupTree.scala 24:34]
  wire [63:0] _T_101 = _T_96 ? msip : 64'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_102 = _T_97 ? freq : 16'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_103 = _T_98 ? mtime : 64'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_104 = _T_99 ? inc : 16'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_105 = _T_100 ? mtimecmp : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _GEN_16 = {{48'd0}, _T_102}; // @[Mux.scala 27:72]
  wire [63:0] _T_106 = _T_101 | _GEN_16; // @[Mux.scala 27:72]
  wire [63:0] _T_107 = _T_106 | _T_103; // @[Mux.scala 27:72]
  wire [63:0] _GEN_17 = {{48'd0}, _T_104}; // @[Mux.scala 27:72]
  wire [63:0] _T_108 = _T_107 | _GEN_17; // @[Mux.scala 27:72]
  wire  _T_111 = io__in_aw_bits_addr[15:0] == 16'h0; // @[RegMap.scala 32:41]
  wire  _T_112 = _T_50 & _T_111; // @[RegMap.scala 32:32]
  wire [63:0] _T_113 = io__in_w_bits_data & fullMask; // @[BitUtils.scala 32:13]
  wire [63:0] _T_114 = ~fullMask; // @[BitUtils.scala 32:38]
  wire [63:0] _T_115 = msip & _T_114; // @[BitUtils.scala 32:36]
  wire [63:0] _T_116 = _T_113 | _T_115; // @[BitUtils.scala 32:25]
  wire  _T_117 = io__in_aw_bits_addr[15:0] == 16'h8000; // @[RegMap.scala 32:41]
  wire  _T_118 = _T_50 & _T_117; // @[RegMap.scala 32:32]
  wire [63:0] _GEN_18 = {{48'd0}, freq}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_121 = _GEN_18 & _T_114; // @[BitUtils.scala 32:36]
  wire [63:0] _T_122 = _T_113 | _T_121; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_11 = _T_118 ? _T_122 : {{48'd0}, freq}; // @[RegMap.scala 32:48]
  wire  _T_123 = io__in_aw_bits_addr[15:0] == 16'hbff8; // @[RegMap.scala 32:41]
  wire  _T_124 = _T_50 & _T_123; // @[RegMap.scala 32:32]
  wire [63:0] _T_127 = mtime & _T_114; // @[BitUtils.scala 32:36]
  wire [63:0] _T_128 = _T_113 | _T_127; // @[BitUtils.scala 32:25]
  wire  _T_129 = io__in_aw_bits_addr[15:0] == 16'h8008; // @[RegMap.scala 32:41]
  wire  _T_130 = _T_50 & _T_129; // @[RegMap.scala 32:32]
  wire [63:0] _T_133 = _GEN_15 & _T_114; // @[BitUtils.scala 32:36]
  wire [63:0] _T_134 = _T_113 | _T_133; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_13 = _T_130 ? _T_134 : {{48'd0}, inc}; // @[RegMap.scala 32:48]
  wire  _T_135 = io__in_aw_bits_addr[15:0] == 16'h4000; // @[RegMap.scala 32:41]
  wire  _T_136 = _T_50 & _T_135; // @[RegMap.scala 32:32]
  wire [63:0] _T_139 = mtimecmp & _T_114; // @[BitUtils.scala 32:36]
  wire [63:0] _T_140 = _T_113 | _T_139; // @[BitUtils.scala 32:25]
  reg  _T_142; // @[AXI4CLINT.scala 64:31]
  reg  _T_144; // @[AXI4CLINT.scala 65:31]
  assign io__in_aw_ready = ~w_busy; // @[AXI4Slave.scala 94:15]
  assign io__in_w_ready = io__in_aw_valid | w_busy; // @[AXI4Slave.scala 95:15]
  assign io__in_b_valid = _T_53; // @[AXI4Slave.scala 97:14]
  assign io__in_ar_ready = io__in_r_ready | _T_33; // @[AXI4Slave.scala 71:15]
  assign io__in_r_valid = _T_45; // @[AXI4Slave.scala 74:14]
  assign io__in_r_bits_data = _T_108 | _T_105; // @[RegMap.scala 30:11]
  assign io__extra_mtip = _T_142; // @[AXI4CLINT.scala 64:21]
  assign io__extra_msip = _T_144; // @[AXI4CLINT.scala 65:21]
  assign io_extra_mtip = io__extra_mtip;
  assign io_extra_msip = io__extra_msip;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ren = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _T_45 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_53 = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  mtime = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mtimecmp = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  msip = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  freq = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  inc = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  cnt = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  _T_142 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _T_144 = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      r_busy <= 1'h0;
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin
      ren <= 1'h0;
    end else begin
      ren <= _T_30;
    end
    if (reset) begin
      _T_45 <= 1'h0;
    end else begin
      _T_45 <= _GEN_3;
    end
    if (reset) begin
      w_busy <= 1'h0;
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin
      _T_53 <= 1'h0;
    end else begin
      _T_53 <= _GEN_7;
    end
    if (reset) begin
      mtime <= 64'h0;
    end else if (_T_124) begin
      mtime <= _T_128;
    end else if (isWFI) begin
      mtime <= _T_61;
    end else if (tick) begin
      mtime <= _T_58;
    end
    if (reset) begin
      mtimecmp <= 64'h0;
    end else if (_T_136) begin
      mtimecmp <= _T_140;
    end
    if (reset) begin
      msip <= 64'h0;
    end else if (_T_112) begin
      msip <= _T_116;
    end
    if (reset) begin
      freq <= 16'h2710;
    end else begin
      freq <= _GEN_11[15:0];
    end
    if (reset) begin
      inc <= 16'h1;
    end else begin
      inc <= _GEN_13[15:0];
    end
    if (reset) begin
      cnt <= 16'h0;
    end else if (_T_55) begin
      cnt <= nextCnt;
    end else begin
      cnt <= 16'h0;
    end
    _T_142 <= mtime >= mtimecmp;
    _T_144 <= msip != 64'h0;
  end
endmodule
module SimpleBus2AXI4Converter_1(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [3:0]  io_in_req_bits_cmd,
  input  [7:0]  io_in_req_bits_wmask,
  input  [63:0] io_in_req_bits_wdata,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_aw_ready,
  output        io_out_aw_valid,
  output [31:0] io_out_aw_bits_addr,
  input         io_out_w_ready,
  output        io_out_w_valid,
  output [63:0] io_out_w_bits_data,
  output [7:0]  io_out_w_bits_strb,
  output        io_out_b_ready,
  input         io_out_b_valid,
  input         io_out_ar_ready,
  output        io_out_ar_valid,
  output [31:0] io_out_ar_bits_addr,
  output        io_out_r_ready,
  input         io_out_r_valid,
  input  [63:0] io_out_r_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  _T_1 = io_in_req_valid & io_in_req_bits_cmd[1]; // @[ToAXI4.scala 151:38]
  wire  toAXI4Lite = ~_T_1; // @[ToAXI4.scala 151:20]
  wire  _T_5 = toAXI4Lite | reset; // @[ToAXI4.scala 153:9]
  wire  _T_6 = ~_T_5; // @[ToAXI4.scala 153:9]
  wire  _T_8 = io_out_aw_ready & io_out_aw_valid; // @[Decoupled.scala 40:37]
  reg  awAck; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_8 | awAck; // @[StopWatch.scala 30:20]
  wire  _T_12 = io_out_w_ready & io_out_w_valid; // @[Decoupled.scala 40:37]
  wire  _T_13 = _T_8 & _T_12; // @[ToAXI4.scala 189:27]
  reg  wAck; // @[StopWatch.scala 24:20]
  wire  _T_15 = awAck & wAck; // @[ToAXI4.scala 189:63]
  wire  wSend = _T_13 | _T_15; // @[ToAXI4.scala 189:53]
  wire  _GEN_2 = _T_12 | wAck; // @[StopWatch.scala 30:20]
  wire  _T_18 = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 40:37]
  reg  wen; // @[Reg.scala 15:16]
  wire  _T_20 = ~io_in_req_bits_cmd[0]; // @[SimpleBus.scala 73:18]
  wire  _T_22 = ~io_in_req_bits_cmd[3]; // @[SimpleBus.scala 73:29]
  wire  _T_23 = _T_20 & _T_22; // @[SimpleBus.scala 73:26]
  wire  _T_26 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[SimpleBus.scala 103:29]
  wire  _T_27 = ~awAck; // @[ToAXI4.scala 193:36]
  wire  _T_31 = ~wAck; // @[ToAXI4.scala 194:36]
  wire  _T_35 = _T_31 & io_out_w_ready; // @[ToAXI4.scala 195:55]
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _T_35 : io_out_ar_ready; // @[ToAXI4.scala 195:18]
  assign io_in_resp_valid = wen ? io_out_b_valid : io_out_r_valid; // @[ToAXI4.scala 199:19]
  assign io_in_resp_bits_rdata = io_out_r_bits_data; // @[ToAXI4.scala 183:23]
  assign io_out_aw_valid = _T_26 & _T_27; // @[ToAXI4.scala 193:16]
  assign io_out_aw_bits_addr = io_out_ar_bits_addr; // @[ToAXI4.scala 182:6]
  assign io_out_w_valid = _T_26 & _T_31; // @[ToAXI4.scala 194:16]
  assign io_out_w_bits_data = io_in_req_bits_wdata; // @[ToAXI4.scala 160:10]
  assign io_out_w_bits_strb = io_in_req_bits_wmask; // @[ToAXI4.scala 161:10]
  assign io_out_b_ready = io_in_resp_ready; // @[ToAXI4.scala 198:16]
  assign io_out_ar_valid = io_in_req_valid & _T_23; // @[ToAXI4.scala 192:16]
  assign io_out_ar_bits_addr = io_in_req_bits_addr; // @[ToAXI4.scala 158:12]
  assign io_out_r_ready = io_in_resp_ready; // @[ToAXI4.scala 197:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  awAck = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wAck = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wen = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      awAck <= 1'h0;
    end else if (wSend) begin
      awAck <= 1'h0;
    end else begin
      awAck <= _GEN_0;
    end
    if (reset) begin
      wAck <= 1'h0;
    end else if (wSend) begin
      wAck <= 1'h0;
    end else begin
      wAck <= _GEN_2;
    end
    if (_T_18) begin
      wen <= io_in_req_bits_cmd[0];
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:153 assert(toAXI4Lite || toAXI4)\n"); // @[ToAXI4.scala 153:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6) begin
          $fatal; // @[ToAXI4.scala 153:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module AXI4PLIC(
  input         clock,
  input         reset,
  output        io__in_aw_ready,
  input         io__in_aw_valid,
  input  [31:0] io__in_aw_bits_addr,
  output        io__in_w_ready,
  input         io__in_w_valid,
  input  [63:0] io__in_w_bits_data,
  input  [7:0]  io__in_w_bits_strb,
  input         io__in_b_ready,
  output        io__in_b_valid,
  output        io__in_ar_ready,
  input         io__in_ar_valid,
  input  [31:0] io__in_ar_bits_addr,
  input         io__in_r_ready,
  output        io__in_r_valid,
  output [63:0] io__in_r_bits_data,
  input         io__extra_intrVec,
  output        io__extra_meip_0,
  output        io_extra_meip_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire  _T_30 = io__in_ar_ready & io__in_ar_valid; // @[Decoupled.scala 40:37]
  wire  _T_31 = io__in_r_ready & io__in_r_valid; // @[Decoupled.scala 40:37]
  reg  r_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_31 ? 1'h0 : r_busy; // @[StopWatch.scala 26:19]
  wire  _GEN_1 = _T_30 | _GEN_0; // @[StopWatch.scala 27:20]
  wire  _T_33 = ~r_busy; // @[AXI4Slave.scala 71:32]
  reg  ren; // @[AXI4Slave.scala 73:17]
  wire  _T_42 = _T_30 | r_busy; // @[AXI4Slave.scala 74:52]
  wire  _T_43 = ren & _T_42; // @[AXI4Slave.scala 74:35]
  reg  _T_45; // @[StopWatch.scala 24:20]
  wire  _GEN_2 = _T_31 ? 1'h0 : _T_45; // @[StopWatch.scala 26:19]
  wire  _GEN_3 = _T_43 | _GEN_2; // @[StopWatch.scala 27:20]
  wire  _T_46 = io__in_aw_ready & io__in_aw_valid; // @[Decoupled.scala 40:37]
  wire  _T_47 = io__in_b_ready & io__in_b_valid; // @[Decoupled.scala 40:37]
  reg  w_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_4 = _T_47 ? 1'h0 : w_busy; // @[StopWatch.scala 26:19]
  wire  _GEN_5 = _T_46 | _GEN_4; // @[StopWatch.scala 27:20]
  wire  _T_50 = io__in_w_ready & io__in_w_valid; // @[Decoupled.scala 40:37]
  reg  _T_53; // @[StopWatch.scala 24:20]
  wire  _GEN_6 = _T_47 ? 1'h0 : _T_53; // @[StopWatch.scala 26:19]
  wire  _GEN_7 = _T_50 | _GEN_6; // @[StopWatch.scala 27:20]
  reg [31:0] priority_0; // @[AXI4PLIC.scala 37:39]
  reg  pending_0_1; // @[AXI4PLIC.scala 43:46]
  wire [31:0] _T_85 = {16'h0,8'h0,4'h0,2'h0,pending_0_1,1'h0}; // @[Cat.scala 29:58]
  reg [31:0] enable_0_0; // @[AXI4PLIC.scala 48:64]
  reg [31:0] threshold_0; // @[AXI4PLIC.scala 53:40]
  reg  inHandle_1; // @[AXI4PLIC.scala 58:25]
  reg [31:0] claimCompletion_0; // @[AXI4PLIC.scala 64:46]
  wire  _T_89 = io__in_ar_bits_addr[25:0] == 26'h200004; // @[AXI4PLIC.scala 68:46]
  wire  _T_90 = _T_31 & _T_89; // @[AXI4PLIC.scala 68:25]
  wire  _GEN_9 = claimCompletion_0[0] | inHandle_1; // @[AXI4PLIC.scala 68:73]
  wire  _GEN_12 = io__extra_intrVec | pending_0_1; // @[AXI4PLIC.scala 75:17]
  wire [31:0] _T_123 = _T_85 & enable_0_0; // @[AXI4PLIC.scala 81:31]
  wire  _T_124 = _T_123 == 32'h0; // @[AXI4PLIC.scala 82:23]
  wire [4:0] _T_157 = _T_123[30] ? 5'h1e : 5'h1f; // @[Mux.scala 47:69]
  wire [4:0] _T_158 = _T_123[29] ? 5'h1d : _T_157; // @[Mux.scala 47:69]
  wire [4:0] _T_159 = _T_123[28] ? 5'h1c : _T_158; // @[Mux.scala 47:69]
  wire [4:0] _T_160 = _T_123[27] ? 5'h1b : _T_159; // @[Mux.scala 47:69]
  wire [4:0] _T_161 = _T_123[26] ? 5'h1a : _T_160; // @[Mux.scala 47:69]
  wire [4:0] _T_162 = _T_123[25] ? 5'h19 : _T_161; // @[Mux.scala 47:69]
  wire [4:0] _T_163 = _T_123[24] ? 5'h18 : _T_162; // @[Mux.scala 47:69]
  wire [4:0] _T_164 = _T_123[23] ? 5'h17 : _T_163; // @[Mux.scala 47:69]
  wire [4:0] _T_165 = _T_123[22] ? 5'h16 : _T_164; // @[Mux.scala 47:69]
  wire [4:0] _T_166 = _T_123[21] ? 5'h15 : _T_165; // @[Mux.scala 47:69]
  wire [4:0] _T_167 = _T_123[20] ? 5'h14 : _T_166; // @[Mux.scala 47:69]
  wire [4:0] _T_168 = _T_123[19] ? 5'h13 : _T_167; // @[Mux.scala 47:69]
  wire [4:0] _T_169 = _T_123[18] ? 5'h12 : _T_168; // @[Mux.scala 47:69]
  wire [4:0] _T_170 = _T_123[17] ? 5'h11 : _T_169; // @[Mux.scala 47:69]
  wire [4:0] _T_171 = _T_123[16] ? 5'h10 : _T_170; // @[Mux.scala 47:69]
  wire [4:0] _T_172 = _T_123[15] ? 5'hf : _T_171; // @[Mux.scala 47:69]
  wire [4:0] _T_173 = _T_123[14] ? 5'he : _T_172; // @[Mux.scala 47:69]
  wire [4:0] _T_174 = _T_123[13] ? 5'hd : _T_173; // @[Mux.scala 47:69]
  wire [4:0] _T_175 = _T_123[12] ? 5'hc : _T_174; // @[Mux.scala 47:69]
  wire [4:0] _T_176 = _T_123[11] ? 5'hb : _T_175; // @[Mux.scala 47:69]
  wire [4:0] _T_177 = _T_123[10] ? 5'ha : _T_176; // @[Mux.scala 47:69]
  wire [4:0] _T_178 = _T_123[9] ? 5'h9 : _T_177; // @[Mux.scala 47:69]
  wire [4:0] _T_179 = _T_123[8] ? 5'h8 : _T_178; // @[Mux.scala 47:69]
  wire [4:0] _T_180 = _T_123[7] ? 5'h7 : _T_179; // @[Mux.scala 47:69]
  wire [4:0] _T_181 = _T_123[6] ? 5'h6 : _T_180; // @[Mux.scala 47:69]
  wire [4:0] _T_182 = _T_123[5] ? 5'h5 : _T_181; // @[Mux.scala 47:69]
  wire [4:0] _T_183 = _T_123[4] ? 5'h4 : _T_182; // @[Mux.scala 47:69]
  wire [4:0] _T_184 = _T_123[3] ? 5'h3 : _T_183; // @[Mux.scala 47:69]
  wire [4:0] _T_185 = _T_123[2] ? 5'h2 : _T_184; // @[Mux.scala 47:69]
  wire [4:0] _T_186 = _T_123[1] ? 5'h1 : _T_185; // @[Mux.scala 47:69]
  wire [4:0] _T_187 = _T_123[0] ? 5'h0 : _T_186; // @[Mux.scala 47:69]
  wire [4:0] _T_188 = _T_124 ? 5'h0 : _T_187; // @[AXI4PLIC.scala 82:13]
  wire [7:0] _T_193 = io__in_w_bits_strb >> io__in_aw_bits_addr[2:0]; // @[AXI4PLIC.scala 89:78]
  wire [7:0] _T_203 = _T_193[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_205 = _T_193[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_207 = _T_193[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_209 = _T_193[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_211 = _T_193[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_213 = _T_193[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_215 = _T_193[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_217 = _T_193[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_224 = {_T_217,_T_215,_T_213,_T_211,_T_209,_T_207,_T_205,_T_203}; // @[Cat.scala 29:58]
  wire  _T_225 = 26'h1000 == io__in_ar_bits_addr[25:0]; // @[LookupTree.scala 24:34]
  wire  _T_226 = 26'h2000 == io__in_ar_bits_addr[25:0]; // @[LookupTree.scala 24:34]
  wire  _T_227 = 26'h200004 == io__in_ar_bits_addr[25:0]; // @[LookupTree.scala 24:34]
  wire  _T_228 = 26'h4 == io__in_ar_bits_addr[25:0]; // @[LookupTree.scala 24:34]
  wire  _T_229 = 26'h200000 == io__in_ar_bits_addr[25:0]; // @[LookupTree.scala 24:34]
  wire [31:0] _T_230 = _T_225 ? _T_85 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_231 = _T_226 ? enable_0_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_232 = _T_227 ? claimCompletion_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_233 = _T_228 ? priority_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_234 = _T_229 ? threshold_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_235 = _T_230 | _T_231; // @[Mux.scala 27:72]
  wire [31:0] _T_236 = _T_235 | _T_232; // @[Mux.scala 27:72]
  wire [31:0] _T_237 = _T_236 | _T_233; // @[Mux.scala 27:72]
  wire [31:0] rdata = _T_237 | _T_234; // @[Mux.scala 27:72]
  wire  _T_240 = io__in_aw_bits_addr[25:0] == 26'h2000; // @[RegMap.scala 32:41]
  wire  _T_241 = _T_50 & _T_240; // @[RegMap.scala 32:32]
  wire [63:0] _T_242 = io__in_w_bits_data & _T_224; // @[BitUtils.scala 32:13]
  wire [63:0] _T_243 = ~_T_224; // @[BitUtils.scala 32:38]
  wire [63:0] _GEN_23 = {{32'd0}, enable_0_0}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_244 = _GEN_23 & _T_243; // @[BitUtils.scala 32:36]
  wire [63:0] _T_245 = _T_242 | _T_244; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_14 = _T_241 ? _T_245 : {{32'd0}, enable_0_0}; // @[RegMap.scala 32:48]
  wire  _T_246 = io__in_aw_bits_addr[25:0] == 26'h200004; // @[RegMap.scala 32:41]
  wire  _T_247 = _T_50 & _T_246; // @[RegMap.scala 32:32]
  wire [63:0] _GEN_24 = {{32'd0}, claimCompletion_0}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_250 = _GEN_24 & _T_243; // @[BitUtils.scala 32:36]
  wire [63:0] _T_251 = _T_242 | _T_250; // @[BitUtils.scala 32:25]
  wire [4:0] _GEN_19 = _T_247 ? 5'h0 : _T_188; // @[RegMap.scala 32:48]
  wire  _T_254 = io__in_aw_bits_addr[25:0] == 26'h4; // @[RegMap.scala 32:41]
  wire  _T_255 = _T_50 & _T_254; // @[RegMap.scala 32:32]
  wire [63:0] _GEN_25 = {{32'd0}, priority_0}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_258 = _GEN_25 & _T_243; // @[BitUtils.scala 32:36]
  wire [63:0] _T_259 = _T_242 | _T_258; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_20 = _T_255 ? _T_259 : {{32'd0}, priority_0}; // @[RegMap.scala 32:48]
  wire  _T_260 = io__in_aw_bits_addr[25:0] == 26'h200000; // @[RegMap.scala 32:41]
  wire  _T_261 = _T_50 & _T_260; // @[RegMap.scala 32:32]
  wire [63:0] _GEN_26 = {{32'd0}, threshold_0}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_264 = _GEN_26 & _T_243; // @[BitUtils.scala 32:36]
  wire [63:0] _T_265 = _T_242 | _T_264; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_21 = _T_261 ? _T_265 : {{32'd0}, threshold_0}; // @[RegMap.scala 32:48]
  assign io__in_aw_ready = ~w_busy; // @[AXI4Slave.scala 94:15]
  assign io__in_w_ready = io__in_aw_valid | w_busy; // @[AXI4Slave.scala 95:15]
  assign io__in_b_valid = _T_53; // @[AXI4Slave.scala 97:14]
  assign io__in_ar_ready = io__in_r_ready | _T_33; // @[AXI4Slave.scala 71:15]
  assign io__in_r_valid = _T_45; // @[AXI4Slave.scala 74:14]
  assign io__in_r_bits_data = {rdata,rdata}; // @[AXI4PLIC.scala 91:18]
  assign io__extra_meip_0 = claimCompletion_0 != 32'h0; // @[AXI4PLIC.scala 93:62]
  assign io_extra_meip_0 = io__extra_meip_0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ren = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _T_45 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_53 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  priority_0 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  pending_0_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  enable_0_0 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  threshold_0 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  inHandle_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  claimCompletion_0 = _RAND_10[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      r_busy <= 1'h0;
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin
      ren <= 1'h0;
    end else begin
      ren <= _T_30;
    end
    if (reset) begin
      _T_45 <= 1'h0;
    end else begin
      _T_45 <= _GEN_3;
    end
    if (reset) begin
      w_busy <= 1'h0;
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin
      _T_53 <= 1'h0;
    end else begin
      _T_53 <= _GEN_7;
    end
    priority_0 <= _GEN_20[31:0];
    if (reset) begin
      pending_0_1 <= 1'h0;
    end else if (inHandle_1) begin
      pending_0_1 <= 1'h0;
    end else begin
      pending_0_1 <= _GEN_12;
    end
    if (reset) begin
      enable_0_0 <= 32'h0;
    end else begin
      enable_0_0 <= _GEN_14[31:0];
    end
    threshold_0 <= _GEN_21[31:0];
    if (reset) begin
      inHandle_1 <= 1'h0;
    end else if (_T_247) begin
      if (_T_251[0]) begin
        inHandle_1 <= 1'h0;
      end else if (_T_90) begin
        inHandle_1 <= _GEN_9;
      end
    end else if (_T_90) begin
      inHandle_1 <= _GEN_9;
    end
    claimCompletion_0 <= {{27'd0}, _GEN_19};
  end
endmodule
module NutShell(
  input         clock,
  input         reset,
  input         io_mem_aw_ready,
  output        io_mem_aw_valid,
  output [31:0] io_mem_aw_bits_addr,
  output [7:0]  io_mem_aw_bits_len,
  output [2:0]  io_mem_aw_bits_size,
  output [1:0]  io_mem_aw_bits_burst,
  input         io_mem_w_ready,
  output        io_mem_w_valid,
  output [63:0] io_mem_w_bits_data,
  output        io_mem_w_bits_last,
  input         io_mem_b_valid,
  input         io_mem_ar_ready,
  output        io_mem_ar_valid,
  output [31:0] io_mem_ar_bits_addr,
  output [7:0]  io_mem_ar_bits_len,
  input         io_mem_r_valid,
  input  [63:0] io_mem_r_bits_data,
  input         io_mem_r_bits_last,
  input         io_mmio_req_ready,
  output        io_mmio_req_valid,
  output [31:0] io_mmio_req_bits_addr,
  output [2:0]  io_mmio_req_bits_size,
  output [3:0]  io_mmio_req_bits_cmd,
  output [7:0]  io_mmio_req_bits_wmask,
  output [63:0] io_mmio_req_bits_wdata,
  output        io_mmio_resp_ready,
  input         io_mmio_resp_valid,
  input  [63:0] io_mmio_resp_bits_rdata,
  output        io_frontend_aw_ready,
  input         io_frontend_aw_valid,
  input  [31:0] io_frontend_aw_bits_addr,
  input  [7:0]  io_frontend_aw_bits_len,
  input  [2:0]  io_frontend_aw_bits_size,
  output        io_frontend_w_ready,
  input         io_frontend_w_valid,
  input  [63:0] io_frontend_w_bits_data,
  input  [7:0]  io_frontend_w_bits_strb,
  input         io_frontend_b_ready,
  output        io_frontend_b_valid,
  output        io_frontend_ar_ready,
  input         io_frontend_ar_valid,
  input  [31:0] io_frontend_ar_bits_addr,
  input         io_frontend_r_ready,
  output        io_frontend_r_valid,
  output [63:0] io_frontend_r_bits_data,
  input         io_meip,
  output [63:0] _T_4181,
  output [63:0] _T_4184,
  output [63:0] _T_4185,
  output        falseWire,
  output        falseWire_0,
  output [1:0]  _T_4178,
  output [63:0] _T_284_0,
  output [63:0] _T_284_1,
  output [63:0] _T_284_2,
  output [63:0] _T_284_3,
  output [63:0] _T_284_4,
  output [63:0] _T_284_5,
  output [63:0] _T_284_6,
  output [63:0] _T_284_7,
  output [63:0] _T_284_8,
  output [63:0] _T_284_9,
  output [63:0] _T_284_10,
  output [63:0] _T_284_11,
  output [63:0] _T_284_12,
  output [63:0] _T_284_13,
  output [63:0] _T_284_14,
  output [63:0] _T_284_15,
  output [63:0] _T_284_16,
  output [63:0] _T_284_17,
  output [63:0] _T_284_18,
  output [63:0] _T_284_19,
  output [63:0] _T_284_20,
  output [63:0] _T_284_21,
  output [63:0] _T_284_22,
  output [63:0] _T_284_23,
  output [63:0] _T_284_24,
  output [63:0] _T_284_25,
  output [63:0] _T_284_26,
  output [63:0] _T_284_27,
  output [63:0] _T_284_28,
  output [63:0] _T_284_29,
  output [63:0] _T_284_30,
  output [63:0] _T_284_31,
  output        _T_36,
  output [63:0] _T_32,
  input         _T_13,
  output [63:0] _T_31,
  output [63:0] _T_37,
  output        _T_26,
  output [63:0] _T_4183,
  output [63:0] _T_4182,
  output        _T_33,
  output [63:0] _T_4179
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  nutcore_clock; // @[NutShell.scala 53:23]
  wire  nutcore_reset; // @[NutShell.scala 53:23]
  wire  nutcore_io_imem_mem_req_ready; // @[NutShell.scala 53:23]
  wire  nutcore_io_imem_mem_req_valid; // @[NutShell.scala 53:23]
  wire [31:0] nutcore_io_imem_mem_req_bits_addr; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_imem_mem_req_bits_cmd; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_imem_mem_req_bits_wdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_imem_mem_resp_valid; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_imem_mem_resp_bits_cmd; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_imem_mem_resp_bits_rdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_dmem_mem_req_ready; // @[NutShell.scala 53:23]
  wire  nutcore_io_dmem_mem_req_valid; // @[NutShell.scala 53:23]
  wire [31:0] nutcore_io_dmem_mem_req_bits_addr; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_dmem_mem_req_bits_cmd; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_dmem_mem_req_bits_wdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_dmem_mem_resp_valid; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_dmem_mem_resp_bits_cmd; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_dmem_mem_resp_bits_rdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_dmem_coh_req_ready; // @[NutShell.scala 53:23]
  wire  nutcore_io_dmem_coh_req_valid; // @[NutShell.scala 53:23]
  wire [31:0] nutcore_io_dmem_coh_req_bits_addr; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_dmem_coh_req_bits_wdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_dmem_coh_resp_valid; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_dmem_coh_resp_bits_cmd; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_dmem_coh_resp_bits_rdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_mmio_req_ready; // @[NutShell.scala 53:23]
  wire  nutcore_io_mmio_req_valid; // @[NutShell.scala 53:23]
  wire [31:0] nutcore_io_mmio_req_bits_addr; // @[NutShell.scala 53:23]
  wire [2:0] nutcore_io_mmio_req_bits_size; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_mmio_req_bits_cmd; // @[NutShell.scala 53:23]
  wire [7:0] nutcore_io_mmio_req_bits_wmask; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_mmio_req_bits_wdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_mmio_resp_valid; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_mmio_resp_bits_rdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_frontend_req_ready; // @[NutShell.scala 53:23]
  wire  nutcore_io_frontend_req_valid; // @[NutShell.scala 53:23]
  wire [31:0] nutcore_io_frontend_req_bits_addr; // @[NutShell.scala 53:23]
  wire [2:0] nutcore_io_frontend_req_bits_size; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_frontend_req_bits_cmd; // @[NutShell.scala 53:23]
  wire [7:0] nutcore_io_frontend_req_bits_wmask; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_frontend_req_bits_wdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_frontend_resp_ready; // @[NutShell.scala 53:23]
  wire  nutcore_io_frontend_resp_valid; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_frontend_resp_bits_cmd; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_frontend_resp_bits_rdata; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_4181; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_4184; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_4185; // @[NutShell.scala 53:23]
  wire  nutcore_falseWire; // @[NutShell.scala 53:23]
  wire  nutcore_falseWire_0; // @[NutShell.scala 53:23]
  wire [1:0] nutcore__T_4178; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_284_0; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_284_1; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_284_2; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_284_3; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_284_4; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_284_5; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_284_6; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_284_7; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_284_8; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_284_9; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_284_10; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_284_11; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_284_12; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_284_13; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_284_14; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_284_15; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_284_16; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_284_17; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_284_18; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_284_19; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_284_20; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_284_21; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_284_22; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_284_23; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_284_24; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_284_25; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_284_26; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_284_27; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_284_28; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_284_29; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_284_30; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_284_31; // @[NutShell.scala 53:23]
  wire  nutcore__T_36_0; // @[NutShell.scala 53:23]
  wire  nutcore_io_extra_mtip; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_32_0; // @[NutShell.scala 53:23]
  wire  nutcore_DISPLAY_ENABLE; // @[NutShell.scala 53:23]
  wire  nutcore_io_extra_meip_0; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_31_0; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_37_0; // @[NutShell.scala 53:23]
  wire  nutcore__T_26_0; // @[NutShell.scala 53:23]
  wire  nutcore__T_0; // @[NutShell.scala 53:23]
  wire  nutcore_io_extra_msip; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_4183; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_4182; // @[NutShell.scala 53:23]
  wire  nutcore__T_33_0; // @[NutShell.scala 53:23]
  wire [63:0] nutcore__T_4179; // @[NutShell.scala 53:23]
  wire  cohMg_clock; // @[NutShell.scala 54:21]
  wire  cohMg_reset; // @[NutShell.scala 54:21]
  wire  cohMg_io_in_req_ready; // @[NutShell.scala 54:21]
  wire  cohMg_io_in_req_valid; // @[NutShell.scala 54:21]
  wire [31:0] cohMg_io_in_req_bits_addr; // @[NutShell.scala 54:21]
  wire [3:0] cohMg_io_in_req_bits_cmd; // @[NutShell.scala 54:21]
  wire [63:0] cohMg_io_in_req_bits_wdata; // @[NutShell.scala 54:21]
  wire  cohMg_io_in_resp_valid; // @[NutShell.scala 54:21]
  wire [3:0] cohMg_io_in_resp_bits_cmd; // @[NutShell.scala 54:21]
  wire [63:0] cohMg_io_in_resp_bits_rdata; // @[NutShell.scala 54:21]
  wire  cohMg_io_out_mem_req_ready; // @[NutShell.scala 54:21]
  wire  cohMg_io_out_mem_req_valid; // @[NutShell.scala 54:21]
  wire [31:0] cohMg_io_out_mem_req_bits_addr; // @[NutShell.scala 54:21]
  wire [3:0] cohMg_io_out_mem_req_bits_cmd; // @[NutShell.scala 54:21]
  wire [63:0] cohMg_io_out_mem_req_bits_wdata; // @[NutShell.scala 54:21]
  wire  cohMg_io_out_mem_resp_ready; // @[NutShell.scala 54:21]
  wire  cohMg_io_out_mem_resp_valid; // @[NutShell.scala 54:21]
  wire [3:0] cohMg_io_out_mem_resp_bits_cmd; // @[NutShell.scala 54:21]
  wire [63:0] cohMg_io_out_mem_resp_bits_rdata; // @[NutShell.scala 54:21]
  wire  cohMg_io_out_coh_req_ready; // @[NutShell.scala 54:21]
  wire  cohMg_io_out_coh_req_valid; // @[NutShell.scala 54:21]
  wire [31:0] cohMg_io_out_coh_req_bits_addr; // @[NutShell.scala 54:21]
  wire [63:0] cohMg_io_out_coh_req_bits_wdata; // @[NutShell.scala 54:21]
  wire  cohMg_io_out_coh_resp_ready; // @[NutShell.scala 54:21]
  wire  cohMg_io_out_coh_resp_valid; // @[NutShell.scala 54:21]
  wire [3:0] cohMg_io_out_coh_resp_bits_cmd; // @[NutShell.scala 54:21]
  wire [63:0] cohMg_io_out_coh_resp_bits_rdata; // @[NutShell.scala 54:21]
  wire  xbar_clock; // @[NutShell.scala 55:20]
  wire  xbar_reset; // @[NutShell.scala 55:20]
  wire  xbar_io_in_0_req_ready; // @[NutShell.scala 55:20]
  wire  xbar_io_in_0_req_valid; // @[NutShell.scala 55:20]
  wire [31:0] xbar_io_in_0_req_bits_addr; // @[NutShell.scala 55:20]
  wire [3:0] xbar_io_in_0_req_bits_cmd; // @[NutShell.scala 55:20]
  wire [7:0] xbar_io_in_0_req_bits_wmask; // @[NutShell.scala 55:20]
  wire [63:0] xbar_io_in_0_req_bits_wdata; // @[NutShell.scala 55:20]
  wire  xbar_io_in_0_resp_valid; // @[NutShell.scala 55:20]
  wire [3:0] xbar_io_in_0_resp_bits_cmd; // @[NutShell.scala 55:20]
  wire [63:0] xbar_io_in_0_resp_bits_rdata; // @[NutShell.scala 55:20]
  wire  xbar_io_in_1_req_ready; // @[NutShell.scala 55:20]
  wire  xbar_io_in_1_req_valid; // @[NutShell.scala 55:20]
  wire [31:0] xbar_io_in_1_req_bits_addr; // @[NutShell.scala 55:20]
  wire [2:0] xbar_io_in_1_req_bits_size; // @[NutShell.scala 55:20]
  wire [3:0] xbar_io_in_1_req_bits_cmd; // @[NutShell.scala 55:20]
  wire [7:0] xbar_io_in_1_req_bits_wmask; // @[NutShell.scala 55:20]
  wire [63:0] xbar_io_in_1_req_bits_wdata; // @[NutShell.scala 55:20]
  wire  xbar_io_in_1_resp_valid; // @[NutShell.scala 55:20]
  wire [3:0] xbar_io_in_1_resp_bits_cmd; // @[NutShell.scala 55:20]
  wire [63:0] xbar_io_in_1_resp_bits_rdata; // @[NutShell.scala 55:20]
  wire  xbar_io_out_req_ready; // @[NutShell.scala 55:20]
  wire  xbar_io_out_req_valid; // @[NutShell.scala 55:20]
  wire [31:0] xbar_io_out_req_bits_addr; // @[NutShell.scala 55:20]
  wire [2:0] xbar_io_out_req_bits_size; // @[NutShell.scala 55:20]
  wire [3:0] xbar_io_out_req_bits_cmd; // @[NutShell.scala 55:20]
  wire [7:0] xbar_io_out_req_bits_wmask; // @[NutShell.scala 55:20]
  wire [63:0] xbar_io_out_req_bits_wdata; // @[NutShell.scala 55:20]
  wire  xbar_io_out_resp_ready; // @[NutShell.scala 55:20]
  wire  xbar_io_out_resp_valid; // @[NutShell.scala 55:20]
  wire [3:0] xbar_io_out_resp_bits_cmd; // @[NutShell.scala 55:20]
  wire [63:0] xbar_io_out_resp_bits_rdata; // @[NutShell.scala 55:20]
  wire  axi2sb_clock; // @[NutShell.scala 61:22]
  wire  axi2sb_reset; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_aw_ready; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_aw_valid; // @[NutShell.scala 61:22]
  wire [31:0] axi2sb_io_in_aw_bits_addr; // @[NutShell.scala 61:22]
  wire [7:0] axi2sb_io_in_aw_bits_len; // @[NutShell.scala 61:22]
  wire [2:0] axi2sb_io_in_aw_bits_size; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_w_ready; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_w_valid; // @[NutShell.scala 61:22]
  wire [63:0] axi2sb_io_in_w_bits_data; // @[NutShell.scala 61:22]
  wire [7:0] axi2sb_io_in_w_bits_strb; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_b_ready; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_b_valid; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_ar_ready; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_ar_valid; // @[NutShell.scala 61:22]
  wire [31:0] axi2sb_io_in_ar_bits_addr; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_r_ready; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_r_valid; // @[NutShell.scala 61:22]
  wire [63:0] axi2sb_io_in_r_bits_data; // @[NutShell.scala 61:22]
  wire  axi2sb_io_out_req_ready; // @[NutShell.scala 61:22]
  wire  axi2sb_io_out_req_valid; // @[NutShell.scala 61:22]
  wire [31:0] axi2sb_io_out_req_bits_addr; // @[NutShell.scala 61:22]
  wire [2:0] axi2sb_io_out_req_bits_size; // @[NutShell.scala 61:22]
  wire [3:0] axi2sb_io_out_req_bits_cmd; // @[NutShell.scala 61:22]
  wire [7:0] axi2sb_io_out_req_bits_wmask; // @[NutShell.scala 61:22]
  wire [63:0] axi2sb_io_out_req_bits_wdata; // @[NutShell.scala 61:22]
  wire  axi2sb_io_out_resp_ready; // @[NutShell.scala 61:22]
  wire  axi2sb_io_out_resp_valid; // @[NutShell.scala 61:22]
  wire [3:0] axi2sb_io_out_resp_bits_cmd; // @[NutShell.scala 61:22]
  wire [63:0] axi2sb_io_out_resp_bits_rdata; // @[NutShell.scala 61:22]
  wire  Prefetcher_clock; // @[NutShell.scala 73:30]
  wire  Prefetcher_reset; // @[NutShell.scala 73:30]
  wire  Prefetcher_io_in_ready; // @[NutShell.scala 73:30]
  wire  Prefetcher_io_in_valid; // @[NutShell.scala 73:30]
  wire [31:0] Prefetcher_io_in_bits_addr; // @[NutShell.scala 73:30]
  wire [2:0] Prefetcher_io_in_bits_size; // @[NutShell.scala 73:30]
  wire [3:0] Prefetcher_io_in_bits_cmd; // @[NutShell.scala 73:30]
  wire [7:0] Prefetcher_io_in_bits_wmask; // @[NutShell.scala 73:30]
  wire [63:0] Prefetcher_io_in_bits_wdata; // @[NutShell.scala 73:30]
  wire  Prefetcher_io_out_ready; // @[NutShell.scala 73:30]
  wire  Prefetcher_io_out_valid; // @[NutShell.scala 73:30]
  wire [31:0] Prefetcher_io_out_bits_addr; // @[NutShell.scala 73:30]
  wire [2:0] Prefetcher_io_out_bits_size; // @[NutShell.scala 73:30]
  wire [3:0] Prefetcher_io_out_bits_cmd; // @[NutShell.scala 73:30]
  wire [7:0] Prefetcher_io_out_bits_wmask; // @[NutShell.scala 73:30]
  wire [63:0] Prefetcher_io_out_bits_wdata; // @[NutShell.scala 73:30]
  wire  Prefetcher_DISPLAY_ENABLE; // @[NutShell.scala 73:30]
  wire  Cache_clock; // @[Cache.scala 678:35]
  wire  Cache_reset; // @[Cache.scala 678:35]
  wire  Cache_io_in_req_ready; // @[Cache.scala 678:35]
  wire  Cache_io_in_req_valid; // @[Cache.scala 678:35]
  wire [31:0] Cache_io_in_req_bits_addr; // @[Cache.scala 678:35]
  wire [2:0] Cache_io_in_req_bits_size; // @[Cache.scala 678:35]
  wire [3:0] Cache_io_in_req_bits_cmd; // @[Cache.scala 678:35]
  wire [7:0] Cache_io_in_req_bits_wmask; // @[Cache.scala 678:35]
  wire [63:0] Cache_io_in_req_bits_wdata; // @[Cache.scala 678:35]
  wire  Cache_io_in_resp_valid; // @[Cache.scala 678:35]
  wire [3:0] Cache_io_in_resp_bits_cmd; // @[Cache.scala 678:35]
  wire [63:0] Cache_io_in_resp_bits_rdata; // @[Cache.scala 678:35]
  wire  Cache_io_out_mem_req_ready; // @[Cache.scala 678:35]
  wire  Cache_io_out_mem_req_valid; // @[Cache.scala 678:35]
  wire [31:0] Cache_io_out_mem_req_bits_addr; // @[Cache.scala 678:35]
  wire [3:0] Cache_io_out_mem_req_bits_cmd; // @[Cache.scala 678:35]
  wire [63:0] Cache_io_out_mem_req_bits_wdata; // @[Cache.scala 678:35]
  wire  Cache_io_out_mem_resp_valid; // @[Cache.scala 678:35]
  wire [3:0] Cache_io_out_mem_resp_bits_cmd; // @[Cache.scala 678:35]
  wire [63:0] Cache_io_out_mem_resp_bits_rdata; // @[Cache.scala 678:35]
  wire  Cache_DISPLAY_ENABLE; // @[Cache.scala 678:35]
  wire  memAddrMap_io_in_req_ready; // @[NutShell.scala 93:26]
  wire  memAddrMap_io_in_req_valid; // @[NutShell.scala 93:26]
  wire [31:0] memAddrMap_io_in_req_bits_addr; // @[NutShell.scala 93:26]
  wire [3:0] memAddrMap_io_in_req_bits_cmd; // @[NutShell.scala 93:26]
  wire [63:0] memAddrMap_io_in_req_bits_wdata; // @[NutShell.scala 93:26]
  wire  memAddrMap_io_in_resp_valid; // @[NutShell.scala 93:26]
  wire [3:0] memAddrMap_io_in_resp_bits_cmd; // @[NutShell.scala 93:26]
  wire [63:0] memAddrMap_io_in_resp_bits_rdata; // @[NutShell.scala 93:26]
  wire  memAddrMap_io_out_req_ready; // @[NutShell.scala 93:26]
  wire  memAddrMap_io_out_req_valid; // @[NutShell.scala 93:26]
  wire [31:0] memAddrMap_io_out_req_bits_addr; // @[NutShell.scala 93:26]
  wire [3:0] memAddrMap_io_out_req_bits_cmd; // @[NutShell.scala 93:26]
  wire [63:0] memAddrMap_io_out_req_bits_wdata; // @[NutShell.scala 93:26]
  wire  memAddrMap_io_out_resp_valid; // @[NutShell.scala 93:26]
  wire [3:0] memAddrMap_io_out_resp_bits_cmd; // @[NutShell.scala 93:26]
  wire [63:0] memAddrMap_io_out_resp_bits_rdata; // @[NutShell.scala 93:26]
  wire  SimpleBus2AXI4Converter_clock; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_reset; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_in_req_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_in_req_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_io_in_req_bits_addr; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_io_in_req_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_io_in_req_bits_wdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_in_resp_valid; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_io_in_resp_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_io_in_resp_bits_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_aw_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_aw_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_io_out_aw_bits_addr; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_io_out_aw_bits_len; // @[ToAXI4.scala 204:24]
  wire [2:0] SimpleBus2AXI4Converter_io_out_aw_bits_size; // @[ToAXI4.scala 204:24]
  wire [1:0] SimpleBus2AXI4Converter_io_out_aw_bits_burst; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_w_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_w_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_io_out_w_bits_data; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_w_bits_last; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_b_valid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_ar_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_ar_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_io_out_ar_bits_addr; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_io_out_ar_bits_len; // @[ToAXI4.scala 204:24]
  wire [2:0] SimpleBus2AXI4Converter_io_out_ar_bits_size; // @[ToAXI4.scala 204:24]
  wire [1:0] SimpleBus2AXI4Converter_io_out_ar_bits_burst; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_r_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_io_out_r_bits_data; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_r_bits_last; // @[ToAXI4.scala 204:24]
  wire  mmioXbar_clock; // @[NutShell.scala 106:24]
  wire  mmioXbar_reset; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_in_req_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_in_req_valid; // @[NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_in_req_bits_addr; // @[NutShell.scala 106:24]
  wire [2:0] mmioXbar_io_in_req_bits_size; // @[NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_in_req_bits_cmd; // @[NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_in_req_bits_wmask; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_in_req_bits_wdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_in_resp_valid; // @[NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_in_resp_bits_cmd; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_in_resp_bits_rdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_req_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_req_valid; // @[NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_out_0_req_bits_addr; // @[NutShell.scala 106:24]
  wire [2:0] mmioXbar_io_out_0_req_bits_size; // @[NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_0_req_bits_cmd; // @[NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_out_0_req_bits_wmask; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_0_req_bits_wdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_resp_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_resp_valid; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_0_resp_bits_rdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_req_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_req_valid; // @[NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_out_1_req_bits_addr; // @[NutShell.scala 106:24]
  wire [2:0] mmioXbar_io_out_1_req_bits_size; // @[NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_1_req_bits_cmd; // @[NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_out_1_req_bits_wmask; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_1_req_bits_wdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_resp_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_resp_valid; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_1_resp_bits_rdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_req_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_req_valid; // @[NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_out_2_req_bits_addr; // @[NutShell.scala 106:24]
  wire [2:0] mmioXbar_io_out_2_req_bits_size; // @[NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_2_req_bits_cmd; // @[NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_out_2_req_bits_wmask; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_2_req_bits_wdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_resp_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_resp_valid; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_2_resp_bits_rdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_DISPLAY_ENABLE; // @[NutShell.scala 106:24]
  wire  clint_clock; // @[NutShell.scala 113:21]
  wire  clint_reset; // @[NutShell.scala 113:21]
  wire  clint_io__in_aw_ready; // @[NutShell.scala 113:21]
  wire  clint_io__in_aw_valid; // @[NutShell.scala 113:21]
  wire [31:0] clint_io__in_aw_bits_addr; // @[NutShell.scala 113:21]
  wire  clint_io__in_w_ready; // @[NutShell.scala 113:21]
  wire  clint_io__in_w_valid; // @[NutShell.scala 113:21]
  wire [63:0] clint_io__in_w_bits_data; // @[NutShell.scala 113:21]
  wire [7:0] clint_io__in_w_bits_strb; // @[NutShell.scala 113:21]
  wire  clint_io__in_b_ready; // @[NutShell.scala 113:21]
  wire  clint_io__in_b_valid; // @[NutShell.scala 113:21]
  wire  clint_io__in_ar_ready; // @[NutShell.scala 113:21]
  wire  clint_io__in_ar_valid; // @[NutShell.scala 113:21]
  wire [31:0] clint_io__in_ar_bits_addr; // @[NutShell.scala 113:21]
  wire  clint_io__in_r_ready; // @[NutShell.scala 113:21]
  wire  clint_io__in_r_valid; // @[NutShell.scala 113:21]
  wire [63:0] clint_io__in_r_bits_data; // @[NutShell.scala 113:21]
  wire  clint_io__extra_mtip; // @[NutShell.scala 113:21]
  wire  clint_io__extra_msip; // @[NutShell.scala 113:21]
  wire  clint_io_extra_mtip; // @[NutShell.scala 113:21]
  wire  clint_isWFI; // @[NutShell.scala 113:21]
  wire  clint_io_extra_msip; // @[NutShell.scala 113:21]
  wire  SimpleBus2AXI4Converter_1_clock; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_reset; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_in_req_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_in_req_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_1_io_in_req_bits_addr; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_1_io_in_req_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_1_io_in_req_bits_wmask; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_1_io_in_req_bits_wdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_in_resp_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_in_resp_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_1_io_in_resp_bits_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_aw_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_aw_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_1_io_out_aw_bits_addr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_w_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_w_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_1_io_out_w_bits_data; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_1_io_out_w_bits_strb; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_b_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_b_valid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_ar_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_ar_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_1_io_out_ar_bits_addr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_r_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_r_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_1_io_out_r_bits_data; // @[ToAXI4.scala 204:24]
  wire  plic_clock; // @[NutShell.scala 120:20]
  wire  plic_reset; // @[NutShell.scala 120:20]
  wire  plic_io__in_aw_ready; // @[NutShell.scala 120:20]
  wire  plic_io__in_aw_valid; // @[NutShell.scala 120:20]
  wire [31:0] plic_io__in_aw_bits_addr; // @[NutShell.scala 120:20]
  wire  plic_io__in_w_ready; // @[NutShell.scala 120:20]
  wire  plic_io__in_w_valid; // @[NutShell.scala 120:20]
  wire [63:0] plic_io__in_w_bits_data; // @[NutShell.scala 120:20]
  wire [7:0] plic_io__in_w_bits_strb; // @[NutShell.scala 120:20]
  wire  plic_io__in_b_ready; // @[NutShell.scala 120:20]
  wire  plic_io__in_b_valid; // @[NutShell.scala 120:20]
  wire  plic_io__in_ar_ready; // @[NutShell.scala 120:20]
  wire  plic_io__in_ar_valid; // @[NutShell.scala 120:20]
  wire [31:0] plic_io__in_ar_bits_addr; // @[NutShell.scala 120:20]
  wire  plic_io__in_r_ready; // @[NutShell.scala 120:20]
  wire  plic_io__in_r_valid; // @[NutShell.scala 120:20]
  wire [63:0] plic_io__in_r_bits_data; // @[NutShell.scala 120:20]
  wire  plic_io__extra_intrVec; // @[NutShell.scala 120:20]
  wire  plic_io__extra_meip_0; // @[NutShell.scala 120:20]
  wire  plic_io_extra_meip_0; // @[NutShell.scala 120:20]
  wire  SimpleBus2AXI4Converter_2_clock; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_reset; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_in_req_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_in_req_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_2_io_in_req_bits_addr; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_2_io_in_req_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_2_io_in_req_bits_wmask; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_2_io_in_req_bits_wdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_in_resp_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_in_resp_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_2_io_in_resp_bits_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_aw_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_aw_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_2_io_out_aw_bits_addr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_w_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_w_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_2_io_out_w_bits_data; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_2_io_out_w_bits_strb; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_b_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_b_valid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_ar_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_ar_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_2_io_out_ar_bits_addr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_r_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_r_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_2_io_out_r_bits_data; // @[ToAXI4.scala 204:24]
  reg  _T_4; // @[NutShell.scala 122:47]
  reg  _T_5; // @[NutShell.scala 122:39]
  NutCore nutcore ( // @[NutShell.scala 53:23]
    .clock(nutcore_clock),
    .reset(nutcore_reset),
    .io_imem_mem_req_ready(nutcore_io_imem_mem_req_ready),
    .io_imem_mem_req_valid(nutcore_io_imem_mem_req_valid),
    .io_imem_mem_req_bits_addr(nutcore_io_imem_mem_req_bits_addr),
    .io_imem_mem_req_bits_cmd(nutcore_io_imem_mem_req_bits_cmd),
    .io_imem_mem_req_bits_wdata(nutcore_io_imem_mem_req_bits_wdata),
    .io_imem_mem_resp_valid(nutcore_io_imem_mem_resp_valid),
    .io_imem_mem_resp_bits_cmd(nutcore_io_imem_mem_resp_bits_cmd),
    .io_imem_mem_resp_bits_rdata(nutcore_io_imem_mem_resp_bits_rdata),
    .io_dmem_mem_req_ready(nutcore_io_dmem_mem_req_ready),
    .io_dmem_mem_req_valid(nutcore_io_dmem_mem_req_valid),
    .io_dmem_mem_req_bits_addr(nutcore_io_dmem_mem_req_bits_addr),
    .io_dmem_mem_req_bits_cmd(nutcore_io_dmem_mem_req_bits_cmd),
    .io_dmem_mem_req_bits_wdata(nutcore_io_dmem_mem_req_bits_wdata),
    .io_dmem_mem_resp_valid(nutcore_io_dmem_mem_resp_valid),
    .io_dmem_mem_resp_bits_cmd(nutcore_io_dmem_mem_resp_bits_cmd),
    .io_dmem_mem_resp_bits_rdata(nutcore_io_dmem_mem_resp_bits_rdata),
    .io_dmem_coh_req_ready(nutcore_io_dmem_coh_req_ready),
    .io_dmem_coh_req_valid(nutcore_io_dmem_coh_req_valid),
    .io_dmem_coh_req_bits_addr(nutcore_io_dmem_coh_req_bits_addr),
    .io_dmem_coh_req_bits_wdata(nutcore_io_dmem_coh_req_bits_wdata),
    .io_dmem_coh_resp_valid(nutcore_io_dmem_coh_resp_valid),
    .io_dmem_coh_resp_bits_cmd(nutcore_io_dmem_coh_resp_bits_cmd),
    .io_dmem_coh_resp_bits_rdata(nutcore_io_dmem_coh_resp_bits_rdata),
    .io_mmio_req_ready(nutcore_io_mmio_req_ready),
    .io_mmio_req_valid(nutcore_io_mmio_req_valid),
    .io_mmio_req_bits_addr(nutcore_io_mmio_req_bits_addr),
    .io_mmio_req_bits_size(nutcore_io_mmio_req_bits_size),
    .io_mmio_req_bits_cmd(nutcore_io_mmio_req_bits_cmd),
    .io_mmio_req_bits_wmask(nutcore_io_mmio_req_bits_wmask),
    .io_mmio_req_bits_wdata(nutcore_io_mmio_req_bits_wdata),
    .io_mmio_resp_valid(nutcore_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(nutcore_io_mmio_resp_bits_rdata),
    .io_frontend_req_ready(nutcore_io_frontend_req_ready),
    .io_frontend_req_valid(nutcore_io_frontend_req_valid),
    .io_frontend_req_bits_addr(nutcore_io_frontend_req_bits_addr),
    .io_frontend_req_bits_size(nutcore_io_frontend_req_bits_size),
    .io_frontend_req_bits_cmd(nutcore_io_frontend_req_bits_cmd),
    .io_frontend_req_bits_wmask(nutcore_io_frontend_req_bits_wmask),
    .io_frontend_req_bits_wdata(nutcore_io_frontend_req_bits_wdata),
    .io_frontend_resp_ready(nutcore_io_frontend_resp_ready),
    .io_frontend_resp_valid(nutcore_io_frontend_resp_valid),
    .io_frontend_resp_bits_cmd(nutcore_io_frontend_resp_bits_cmd),
    .io_frontend_resp_bits_rdata(nutcore_io_frontend_resp_bits_rdata),
    ._T_4181(nutcore__T_4181),
    ._T_4184(nutcore__T_4184),
    ._T_4185(nutcore__T_4185),
    .falseWire(nutcore_falseWire),
    .falseWire_0(nutcore_falseWire_0),
    ._T_4178(nutcore__T_4178),
    ._T_284_0(nutcore__T_284_0),
    ._T_284_1(nutcore__T_284_1),
    ._T_284_2(nutcore__T_284_2),
    ._T_284_3(nutcore__T_284_3),
    ._T_284_4(nutcore__T_284_4),
    ._T_284_5(nutcore__T_284_5),
    ._T_284_6(nutcore__T_284_6),
    ._T_284_7(nutcore__T_284_7),
    ._T_284_8(nutcore__T_284_8),
    ._T_284_9(nutcore__T_284_9),
    ._T_284_10(nutcore__T_284_10),
    ._T_284_11(nutcore__T_284_11),
    ._T_284_12(nutcore__T_284_12),
    ._T_284_13(nutcore__T_284_13),
    ._T_284_14(nutcore__T_284_14),
    ._T_284_15(nutcore__T_284_15),
    ._T_284_16(nutcore__T_284_16),
    ._T_284_17(nutcore__T_284_17),
    ._T_284_18(nutcore__T_284_18),
    ._T_284_19(nutcore__T_284_19),
    ._T_284_20(nutcore__T_284_20),
    ._T_284_21(nutcore__T_284_21),
    ._T_284_22(nutcore__T_284_22),
    ._T_284_23(nutcore__T_284_23),
    ._T_284_24(nutcore__T_284_24),
    ._T_284_25(nutcore__T_284_25),
    ._T_284_26(nutcore__T_284_26),
    ._T_284_27(nutcore__T_284_27),
    ._T_284_28(nutcore__T_284_28),
    ._T_284_29(nutcore__T_284_29),
    ._T_284_30(nutcore__T_284_30),
    ._T_284_31(nutcore__T_284_31),
    ._T_36_0(nutcore__T_36_0),
    .io_extra_mtip(nutcore_io_extra_mtip),
    ._T_32_0(nutcore__T_32_0),
    .DISPLAY_ENABLE(nutcore_DISPLAY_ENABLE),
    .io_extra_meip_0(nutcore_io_extra_meip_0),
    ._T_31_0(nutcore__T_31_0),
    ._T_37_0(nutcore__T_37_0),
    ._T_26_0(nutcore__T_26_0),
    ._T_0(nutcore__T_0),
    .io_extra_msip(nutcore_io_extra_msip),
    ._T_4183(nutcore__T_4183),
    ._T_4182(nutcore__T_4182),
    ._T_33_0(nutcore__T_33_0),
    ._T_4179(nutcore__T_4179)
  );
  CoherenceManager cohMg ( // @[NutShell.scala 54:21]
    .clock(cohMg_clock),
    .reset(cohMg_reset),
    .io_in_req_ready(cohMg_io_in_req_ready),
    .io_in_req_valid(cohMg_io_in_req_valid),
    .io_in_req_bits_addr(cohMg_io_in_req_bits_addr),
    .io_in_req_bits_cmd(cohMg_io_in_req_bits_cmd),
    .io_in_req_bits_wdata(cohMg_io_in_req_bits_wdata),
    .io_in_resp_valid(cohMg_io_in_resp_valid),
    .io_in_resp_bits_cmd(cohMg_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(cohMg_io_in_resp_bits_rdata),
    .io_out_mem_req_ready(cohMg_io_out_mem_req_ready),
    .io_out_mem_req_valid(cohMg_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(cohMg_io_out_mem_req_bits_addr),
    .io_out_mem_req_bits_cmd(cohMg_io_out_mem_req_bits_cmd),
    .io_out_mem_req_bits_wdata(cohMg_io_out_mem_req_bits_wdata),
    .io_out_mem_resp_ready(cohMg_io_out_mem_resp_ready),
    .io_out_mem_resp_valid(cohMg_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_cmd(cohMg_io_out_mem_resp_bits_cmd),
    .io_out_mem_resp_bits_rdata(cohMg_io_out_mem_resp_bits_rdata),
    .io_out_coh_req_ready(cohMg_io_out_coh_req_ready),
    .io_out_coh_req_valid(cohMg_io_out_coh_req_valid),
    .io_out_coh_req_bits_addr(cohMg_io_out_coh_req_bits_addr),
    .io_out_coh_req_bits_wdata(cohMg_io_out_coh_req_bits_wdata),
    .io_out_coh_resp_ready(cohMg_io_out_coh_resp_ready),
    .io_out_coh_resp_valid(cohMg_io_out_coh_resp_valid),
    .io_out_coh_resp_bits_cmd(cohMg_io_out_coh_resp_bits_cmd),
    .io_out_coh_resp_bits_rdata(cohMg_io_out_coh_resp_bits_rdata)
  );
  SimpleBusCrossbarNto1 xbar ( // @[NutShell.scala 55:20]
    .clock(xbar_clock),
    .reset(xbar_reset),
    .io_in_0_req_ready(xbar_io_in_0_req_ready),
    .io_in_0_req_valid(xbar_io_in_0_req_valid),
    .io_in_0_req_bits_addr(xbar_io_in_0_req_bits_addr),
    .io_in_0_req_bits_cmd(xbar_io_in_0_req_bits_cmd),
    .io_in_0_req_bits_wmask(xbar_io_in_0_req_bits_wmask),
    .io_in_0_req_bits_wdata(xbar_io_in_0_req_bits_wdata),
    .io_in_0_resp_valid(xbar_io_in_0_resp_valid),
    .io_in_0_resp_bits_cmd(xbar_io_in_0_resp_bits_cmd),
    .io_in_0_resp_bits_rdata(xbar_io_in_0_resp_bits_rdata),
    .io_in_1_req_ready(xbar_io_in_1_req_ready),
    .io_in_1_req_valid(xbar_io_in_1_req_valid),
    .io_in_1_req_bits_addr(xbar_io_in_1_req_bits_addr),
    .io_in_1_req_bits_size(xbar_io_in_1_req_bits_size),
    .io_in_1_req_bits_cmd(xbar_io_in_1_req_bits_cmd),
    .io_in_1_req_bits_wmask(xbar_io_in_1_req_bits_wmask),
    .io_in_1_req_bits_wdata(xbar_io_in_1_req_bits_wdata),
    .io_in_1_resp_valid(xbar_io_in_1_resp_valid),
    .io_in_1_resp_bits_cmd(xbar_io_in_1_resp_bits_cmd),
    .io_in_1_resp_bits_rdata(xbar_io_in_1_resp_bits_rdata),
    .io_out_req_ready(xbar_io_out_req_ready),
    .io_out_req_valid(xbar_io_out_req_valid),
    .io_out_req_bits_addr(xbar_io_out_req_bits_addr),
    .io_out_req_bits_size(xbar_io_out_req_bits_size),
    .io_out_req_bits_cmd(xbar_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(xbar_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(xbar_io_out_req_bits_wdata),
    .io_out_resp_ready(xbar_io_out_resp_ready),
    .io_out_resp_valid(xbar_io_out_resp_valid),
    .io_out_resp_bits_cmd(xbar_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(xbar_io_out_resp_bits_rdata)
  );
  AXI42SimpleBusConverter axi2sb ( // @[NutShell.scala 61:22]
    .clock(axi2sb_clock),
    .reset(axi2sb_reset),
    .io_in_aw_ready(axi2sb_io_in_aw_ready),
    .io_in_aw_valid(axi2sb_io_in_aw_valid),
    .io_in_aw_bits_addr(axi2sb_io_in_aw_bits_addr),
    .io_in_aw_bits_len(axi2sb_io_in_aw_bits_len),
    .io_in_aw_bits_size(axi2sb_io_in_aw_bits_size),
    .io_in_w_ready(axi2sb_io_in_w_ready),
    .io_in_w_valid(axi2sb_io_in_w_valid),
    .io_in_w_bits_data(axi2sb_io_in_w_bits_data),
    .io_in_w_bits_strb(axi2sb_io_in_w_bits_strb),
    .io_in_b_ready(axi2sb_io_in_b_ready),
    .io_in_b_valid(axi2sb_io_in_b_valid),
    .io_in_ar_ready(axi2sb_io_in_ar_ready),
    .io_in_ar_valid(axi2sb_io_in_ar_valid),
    .io_in_ar_bits_addr(axi2sb_io_in_ar_bits_addr),
    .io_in_r_ready(axi2sb_io_in_r_ready),
    .io_in_r_valid(axi2sb_io_in_r_valid),
    .io_in_r_bits_data(axi2sb_io_in_r_bits_data),
    .io_out_req_ready(axi2sb_io_out_req_ready),
    .io_out_req_valid(axi2sb_io_out_req_valid),
    .io_out_req_bits_addr(axi2sb_io_out_req_bits_addr),
    .io_out_req_bits_size(axi2sb_io_out_req_bits_size),
    .io_out_req_bits_cmd(axi2sb_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(axi2sb_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(axi2sb_io_out_req_bits_wdata),
    .io_out_resp_ready(axi2sb_io_out_resp_ready),
    .io_out_resp_valid(axi2sb_io_out_resp_valid),
    .io_out_resp_bits_cmd(axi2sb_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(axi2sb_io_out_resp_bits_rdata)
  );
  Prefetcher Prefetcher ( // @[NutShell.scala 73:30]
    .clock(Prefetcher_clock),
    .reset(Prefetcher_reset),
    .io_in_ready(Prefetcher_io_in_ready),
    .io_in_valid(Prefetcher_io_in_valid),
    .io_in_bits_addr(Prefetcher_io_in_bits_addr),
    .io_in_bits_size(Prefetcher_io_in_bits_size),
    .io_in_bits_cmd(Prefetcher_io_in_bits_cmd),
    .io_in_bits_wmask(Prefetcher_io_in_bits_wmask),
    .io_in_bits_wdata(Prefetcher_io_in_bits_wdata),
    .io_out_ready(Prefetcher_io_out_ready),
    .io_out_valid(Prefetcher_io_out_valid),
    .io_out_bits_addr(Prefetcher_io_out_bits_addr),
    .io_out_bits_size(Prefetcher_io_out_bits_size),
    .io_out_bits_cmd(Prefetcher_io_out_bits_cmd),
    .io_out_bits_wmask(Prefetcher_io_out_bits_wmask),
    .io_out_bits_wdata(Prefetcher_io_out_bits_wdata),
    .DISPLAY_ENABLE(Prefetcher_DISPLAY_ENABLE)
  );
  Cache_2 Cache ( // @[Cache.scala 678:35]
    .clock(Cache_clock),
    .reset(Cache_reset),
    .io_in_req_ready(Cache_io_in_req_ready),
    .io_in_req_valid(Cache_io_in_req_valid),
    .io_in_req_bits_addr(Cache_io_in_req_bits_addr),
    .io_in_req_bits_size(Cache_io_in_req_bits_size),
    .io_in_req_bits_cmd(Cache_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(Cache_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(Cache_io_in_req_bits_wdata),
    .io_in_resp_valid(Cache_io_in_resp_valid),
    .io_in_resp_bits_cmd(Cache_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(Cache_io_in_resp_bits_rdata),
    .io_out_mem_req_ready(Cache_io_out_mem_req_ready),
    .io_out_mem_req_valid(Cache_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(Cache_io_out_mem_req_bits_addr),
    .io_out_mem_req_bits_cmd(Cache_io_out_mem_req_bits_cmd),
    .io_out_mem_req_bits_wdata(Cache_io_out_mem_req_bits_wdata),
    .io_out_mem_resp_valid(Cache_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_cmd(Cache_io_out_mem_resp_bits_cmd),
    .io_out_mem_resp_bits_rdata(Cache_io_out_mem_resp_bits_rdata),
    .DISPLAY_ENABLE(Cache_DISPLAY_ENABLE)
  );
  SimpleBusAddressMapper memAddrMap ( // @[NutShell.scala 93:26]
    .io_in_req_ready(memAddrMap_io_in_req_ready),
    .io_in_req_valid(memAddrMap_io_in_req_valid),
    .io_in_req_bits_addr(memAddrMap_io_in_req_bits_addr),
    .io_in_req_bits_cmd(memAddrMap_io_in_req_bits_cmd),
    .io_in_req_bits_wdata(memAddrMap_io_in_req_bits_wdata),
    .io_in_resp_valid(memAddrMap_io_in_resp_valid),
    .io_in_resp_bits_cmd(memAddrMap_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(memAddrMap_io_in_resp_bits_rdata),
    .io_out_req_ready(memAddrMap_io_out_req_ready),
    .io_out_req_valid(memAddrMap_io_out_req_valid),
    .io_out_req_bits_addr(memAddrMap_io_out_req_bits_addr),
    .io_out_req_bits_cmd(memAddrMap_io_out_req_bits_cmd),
    .io_out_req_bits_wdata(memAddrMap_io_out_req_bits_wdata),
    .io_out_resp_valid(memAddrMap_io_out_resp_valid),
    .io_out_resp_bits_cmd(memAddrMap_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(memAddrMap_io_out_resp_bits_rdata)
  );
  SimpleBus2AXI4Converter SimpleBus2AXI4Converter ( // @[ToAXI4.scala 204:24]
    .clock(SimpleBus2AXI4Converter_clock),
    .reset(SimpleBus2AXI4Converter_reset),
    .io_in_req_ready(SimpleBus2AXI4Converter_io_in_req_ready),
    .io_in_req_valid(SimpleBus2AXI4Converter_io_in_req_valid),
    .io_in_req_bits_addr(SimpleBus2AXI4Converter_io_in_req_bits_addr),
    .io_in_req_bits_cmd(SimpleBus2AXI4Converter_io_in_req_bits_cmd),
    .io_in_req_bits_wdata(SimpleBus2AXI4Converter_io_in_req_bits_wdata),
    .io_in_resp_valid(SimpleBus2AXI4Converter_io_in_resp_valid),
    .io_in_resp_bits_cmd(SimpleBus2AXI4Converter_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(SimpleBus2AXI4Converter_io_in_resp_bits_rdata),
    .io_out_aw_ready(SimpleBus2AXI4Converter_io_out_aw_ready),
    .io_out_aw_valid(SimpleBus2AXI4Converter_io_out_aw_valid),
    .io_out_aw_bits_addr(SimpleBus2AXI4Converter_io_out_aw_bits_addr),
    .io_out_aw_bits_len(SimpleBus2AXI4Converter_io_out_aw_bits_len),
    .io_out_aw_bits_size(SimpleBus2AXI4Converter_io_out_aw_bits_size),
    .io_out_aw_bits_burst(SimpleBus2AXI4Converter_io_out_aw_bits_burst),
    .io_out_w_ready(SimpleBus2AXI4Converter_io_out_w_ready),
    .io_out_w_valid(SimpleBus2AXI4Converter_io_out_w_valid),
    .io_out_w_bits_data(SimpleBus2AXI4Converter_io_out_w_bits_data),
    .io_out_w_bits_last(SimpleBus2AXI4Converter_io_out_w_bits_last),
    .io_out_b_valid(SimpleBus2AXI4Converter_io_out_b_valid),
    .io_out_ar_ready(SimpleBus2AXI4Converter_io_out_ar_ready),
    .io_out_ar_valid(SimpleBus2AXI4Converter_io_out_ar_valid),
    .io_out_ar_bits_addr(SimpleBus2AXI4Converter_io_out_ar_bits_addr),
    .io_out_ar_bits_len(SimpleBus2AXI4Converter_io_out_ar_bits_len),
    .io_out_ar_bits_size(SimpleBus2AXI4Converter_io_out_ar_bits_size),
    .io_out_ar_bits_burst(SimpleBus2AXI4Converter_io_out_ar_bits_burst),
    .io_out_r_valid(SimpleBus2AXI4Converter_io_out_r_valid),
    .io_out_r_bits_data(SimpleBus2AXI4Converter_io_out_r_bits_data),
    .io_out_r_bits_last(SimpleBus2AXI4Converter_io_out_r_bits_last)
  );
  SimpleBusCrossbar1toN mmioXbar ( // @[NutShell.scala 106:24]
    .clock(mmioXbar_clock),
    .reset(mmioXbar_reset),
    .io_in_req_ready(mmioXbar_io_in_req_ready),
    .io_in_req_valid(mmioXbar_io_in_req_valid),
    .io_in_req_bits_addr(mmioXbar_io_in_req_bits_addr),
    .io_in_req_bits_size(mmioXbar_io_in_req_bits_size),
    .io_in_req_bits_cmd(mmioXbar_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(mmioXbar_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(mmioXbar_io_in_req_bits_wdata),
    .io_in_resp_valid(mmioXbar_io_in_resp_valid),
    .io_in_resp_bits_cmd(mmioXbar_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(mmioXbar_io_in_resp_bits_rdata),
    .io_out_0_req_ready(mmioXbar_io_out_0_req_ready),
    .io_out_0_req_valid(mmioXbar_io_out_0_req_valid),
    .io_out_0_req_bits_addr(mmioXbar_io_out_0_req_bits_addr),
    .io_out_0_req_bits_size(mmioXbar_io_out_0_req_bits_size),
    .io_out_0_req_bits_cmd(mmioXbar_io_out_0_req_bits_cmd),
    .io_out_0_req_bits_wmask(mmioXbar_io_out_0_req_bits_wmask),
    .io_out_0_req_bits_wdata(mmioXbar_io_out_0_req_bits_wdata),
    .io_out_0_resp_ready(mmioXbar_io_out_0_resp_ready),
    .io_out_0_resp_valid(mmioXbar_io_out_0_resp_valid),
    .io_out_0_resp_bits_rdata(mmioXbar_io_out_0_resp_bits_rdata),
    .io_out_1_req_ready(mmioXbar_io_out_1_req_ready),
    .io_out_1_req_valid(mmioXbar_io_out_1_req_valid),
    .io_out_1_req_bits_addr(mmioXbar_io_out_1_req_bits_addr),
    .io_out_1_req_bits_size(mmioXbar_io_out_1_req_bits_size),
    .io_out_1_req_bits_cmd(mmioXbar_io_out_1_req_bits_cmd),
    .io_out_1_req_bits_wmask(mmioXbar_io_out_1_req_bits_wmask),
    .io_out_1_req_bits_wdata(mmioXbar_io_out_1_req_bits_wdata),
    .io_out_1_resp_ready(mmioXbar_io_out_1_resp_ready),
    .io_out_1_resp_valid(mmioXbar_io_out_1_resp_valid),
    .io_out_1_resp_bits_rdata(mmioXbar_io_out_1_resp_bits_rdata),
    .io_out_2_req_ready(mmioXbar_io_out_2_req_ready),
    .io_out_2_req_valid(mmioXbar_io_out_2_req_valid),
    .io_out_2_req_bits_addr(mmioXbar_io_out_2_req_bits_addr),
    .io_out_2_req_bits_size(mmioXbar_io_out_2_req_bits_size),
    .io_out_2_req_bits_cmd(mmioXbar_io_out_2_req_bits_cmd),
    .io_out_2_req_bits_wmask(mmioXbar_io_out_2_req_bits_wmask),
    .io_out_2_req_bits_wdata(mmioXbar_io_out_2_req_bits_wdata),
    .io_out_2_resp_ready(mmioXbar_io_out_2_resp_ready),
    .io_out_2_resp_valid(mmioXbar_io_out_2_resp_valid),
    .io_out_2_resp_bits_rdata(mmioXbar_io_out_2_resp_bits_rdata),
    .DISPLAY_ENABLE(mmioXbar_DISPLAY_ENABLE)
  );
  AXI4CLINT clint ( // @[NutShell.scala 113:21]
    .clock(clint_clock),
    .reset(clint_reset),
    .io__in_aw_ready(clint_io__in_aw_ready),
    .io__in_aw_valid(clint_io__in_aw_valid),
    .io__in_aw_bits_addr(clint_io__in_aw_bits_addr),
    .io__in_w_ready(clint_io__in_w_ready),
    .io__in_w_valid(clint_io__in_w_valid),
    .io__in_w_bits_data(clint_io__in_w_bits_data),
    .io__in_w_bits_strb(clint_io__in_w_bits_strb),
    .io__in_b_ready(clint_io__in_b_ready),
    .io__in_b_valid(clint_io__in_b_valid),
    .io__in_ar_ready(clint_io__in_ar_ready),
    .io__in_ar_valid(clint_io__in_ar_valid),
    .io__in_ar_bits_addr(clint_io__in_ar_bits_addr),
    .io__in_r_ready(clint_io__in_r_ready),
    .io__in_r_valid(clint_io__in_r_valid),
    .io__in_r_bits_data(clint_io__in_r_bits_data),
    .io__extra_mtip(clint_io__extra_mtip),
    .io__extra_msip(clint_io__extra_msip),
    .io_extra_mtip(clint_io_extra_mtip),
    .isWFI(clint_isWFI),
    .io_extra_msip(clint_io_extra_msip)
  );
  SimpleBus2AXI4Converter_1 SimpleBus2AXI4Converter_1 ( // @[ToAXI4.scala 204:24]
    .clock(SimpleBus2AXI4Converter_1_clock),
    .reset(SimpleBus2AXI4Converter_1_reset),
    .io_in_req_ready(SimpleBus2AXI4Converter_1_io_in_req_ready),
    .io_in_req_valid(SimpleBus2AXI4Converter_1_io_in_req_valid),
    .io_in_req_bits_addr(SimpleBus2AXI4Converter_1_io_in_req_bits_addr),
    .io_in_req_bits_cmd(SimpleBus2AXI4Converter_1_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(SimpleBus2AXI4Converter_1_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(SimpleBus2AXI4Converter_1_io_in_req_bits_wdata),
    .io_in_resp_ready(SimpleBus2AXI4Converter_1_io_in_resp_ready),
    .io_in_resp_valid(SimpleBus2AXI4Converter_1_io_in_resp_valid),
    .io_in_resp_bits_rdata(SimpleBus2AXI4Converter_1_io_in_resp_bits_rdata),
    .io_out_aw_ready(SimpleBus2AXI4Converter_1_io_out_aw_ready),
    .io_out_aw_valid(SimpleBus2AXI4Converter_1_io_out_aw_valid),
    .io_out_aw_bits_addr(SimpleBus2AXI4Converter_1_io_out_aw_bits_addr),
    .io_out_w_ready(SimpleBus2AXI4Converter_1_io_out_w_ready),
    .io_out_w_valid(SimpleBus2AXI4Converter_1_io_out_w_valid),
    .io_out_w_bits_data(SimpleBus2AXI4Converter_1_io_out_w_bits_data),
    .io_out_w_bits_strb(SimpleBus2AXI4Converter_1_io_out_w_bits_strb),
    .io_out_b_ready(SimpleBus2AXI4Converter_1_io_out_b_ready),
    .io_out_b_valid(SimpleBus2AXI4Converter_1_io_out_b_valid),
    .io_out_ar_ready(SimpleBus2AXI4Converter_1_io_out_ar_ready),
    .io_out_ar_valid(SimpleBus2AXI4Converter_1_io_out_ar_valid),
    .io_out_ar_bits_addr(SimpleBus2AXI4Converter_1_io_out_ar_bits_addr),
    .io_out_r_ready(SimpleBus2AXI4Converter_1_io_out_r_ready),
    .io_out_r_valid(SimpleBus2AXI4Converter_1_io_out_r_valid),
    .io_out_r_bits_data(SimpleBus2AXI4Converter_1_io_out_r_bits_data)
  );
  AXI4PLIC plic ( // @[NutShell.scala 120:20]
    .clock(plic_clock),
    .reset(plic_reset),
    .io__in_aw_ready(plic_io__in_aw_ready),
    .io__in_aw_valid(plic_io__in_aw_valid),
    .io__in_aw_bits_addr(plic_io__in_aw_bits_addr),
    .io__in_w_ready(plic_io__in_w_ready),
    .io__in_w_valid(plic_io__in_w_valid),
    .io__in_w_bits_data(plic_io__in_w_bits_data),
    .io__in_w_bits_strb(plic_io__in_w_bits_strb),
    .io__in_b_ready(plic_io__in_b_ready),
    .io__in_b_valid(plic_io__in_b_valid),
    .io__in_ar_ready(plic_io__in_ar_ready),
    .io__in_ar_valid(plic_io__in_ar_valid),
    .io__in_ar_bits_addr(plic_io__in_ar_bits_addr),
    .io__in_r_ready(plic_io__in_r_ready),
    .io__in_r_valid(plic_io__in_r_valid),
    .io__in_r_bits_data(plic_io__in_r_bits_data),
    .io__extra_intrVec(plic_io__extra_intrVec),
    .io__extra_meip_0(plic_io__extra_meip_0),
    .io_extra_meip_0(plic_io_extra_meip_0)
  );
  SimpleBus2AXI4Converter_1 SimpleBus2AXI4Converter_2 ( // @[ToAXI4.scala 204:24]
    .clock(SimpleBus2AXI4Converter_2_clock),
    .reset(SimpleBus2AXI4Converter_2_reset),
    .io_in_req_ready(SimpleBus2AXI4Converter_2_io_in_req_ready),
    .io_in_req_valid(SimpleBus2AXI4Converter_2_io_in_req_valid),
    .io_in_req_bits_addr(SimpleBus2AXI4Converter_2_io_in_req_bits_addr),
    .io_in_req_bits_cmd(SimpleBus2AXI4Converter_2_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(SimpleBus2AXI4Converter_2_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(SimpleBus2AXI4Converter_2_io_in_req_bits_wdata),
    .io_in_resp_ready(SimpleBus2AXI4Converter_2_io_in_resp_ready),
    .io_in_resp_valid(SimpleBus2AXI4Converter_2_io_in_resp_valid),
    .io_in_resp_bits_rdata(SimpleBus2AXI4Converter_2_io_in_resp_bits_rdata),
    .io_out_aw_ready(SimpleBus2AXI4Converter_2_io_out_aw_ready),
    .io_out_aw_valid(SimpleBus2AXI4Converter_2_io_out_aw_valid),
    .io_out_aw_bits_addr(SimpleBus2AXI4Converter_2_io_out_aw_bits_addr),
    .io_out_w_ready(SimpleBus2AXI4Converter_2_io_out_w_ready),
    .io_out_w_valid(SimpleBus2AXI4Converter_2_io_out_w_valid),
    .io_out_w_bits_data(SimpleBus2AXI4Converter_2_io_out_w_bits_data),
    .io_out_w_bits_strb(SimpleBus2AXI4Converter_2_io_out_w_bits_strb),
    .io_out_b_ready(SimpleBus2AXI4Converter_2_io_out_b_ready),
    .io_out_b_valid(SimpleBus2AXI4Converter_2_io_out_b_valid),
    .io_out_ar_ready(SimpleBus2AXI4Converter_2_io_out_ar_ready),
    .io_out_ar_valid(SimpleBus2AXI4Converter_2_io_out_ar_valid),
    .io_out_ar_bits_addr(SimpleBus2AXI4Converter_2_io_out_ar_bits_addr),
    .io_out_r_ready(SimpleBus2AXI4Converter_2_io_out_r_ready),
    .io_out_r_valid(SimpleBus2AXI4Converter_2_io_out_r_valid),
    .io_out_r_bits_data(SimpleBus2AXI4Converter_2_io_out_r_bits_data)
  );
  assign io_mem_aw_valid = SimpleBus2AXI4Converter_io_out_aw_valid; // @[NutShell.scala 95:10]
  assign io_mem_aw_bits_addr = SimpleBus2AXI4Converter_io_out_aw_bits_addr; // @[NutShell.scala 95:10]
  assign io_mem_aw_bits_len = SimpleBus2AXI4Converter_io_out_aw_bits_len; // @[NutShell.scala 95:10]
  assign io_mem_aw_bits_size = SimpleBus2AXI4Converter_io_out_aw_bits_size; // @[NutShell.scala 95:10]
  assign io_mem_aw_bits_burst = SimpleBus2AXI4Converter_io_out_aw_bits_burst; // @[NutShell.scala 95:10]
  assign io_mem_w_valid = SimpleBus2AXI4Converter_io_out_w_valid; // @[NutShell.scala 95:10]
  assign io_mem_w_bits_data = SimpleBus2AXI4Converter_io_out_w_bits_data; // @[NutShell.scala 95:10]
  assign io_mem_w_bits_last = SimpleBus2AXI4Converter_io_out_w_bits_last; // @[NutShell.scala 95:10]
  assign io_mem_ar_valid = SimpleBus2AXI4Converter_io_out_ar_valid; // @[NutShell.scala 95:10]
  assign io_mem_ar_bits_addr = SimpleBus2AXI4Converter_io_out_ar_bits_addr; // @[NutShell.scala 95:10]
  assign io_mem_ar_bits_len = SimpleBus2AXI4Converter_io_out_ar_bits_len; // @[NutShell.scala 95:10]
  assign io_mmio_req_valid = mmioXbar_io_out_0_req_valid; // @[NutShell.scala 111:18]
  assign io_mmio_req_bits_addr = mmioXbar_io_out_0_req_bits_addr; // @[NutShell.scala 111:18]
  assign io_mmio_req_bits_size = mmioXbar_io_out_0_req_bits_size; // @[NutShell.scala 111:18]
  assign io_mmio_req_bits_cmd = mmioXbar_io_out_0_req_bits_cmd; // @[NutShell.scala 111:18]
  assign io_mmio_req_bits_wmask = mmioXbar_io_out_0_req_bits_wmask; // @[NutShell.scala 111:18]
  assign io_mmio_req_bits_wdata = mmioXbar_io_out_0_req_bits_wdata; // @[NutShell.scala 111:18]
  assign io_mmio_resp_ready = mmioXbar_io_out_0_resp_ready; // @[NutShell.scala 111:18]
  assign io_frontend_aw_ready = axi2sb_io_in_aw_ready; // @[NutShell.scala 62:16]
  assign io_frontend_w_ready = axi2sb_io_in_w_ready; // @[NutShell.scala 62:16]
  assign io_frontend_b_valid = axi2sb_io_in_b_valid; // @[NutShell.scala 62:16]
  assign io_frontend_ar_ready = axi2sb_io_in_ar_ready; // @[NutShell.scala 62:16]
  assign io_frontend_r_valid = axi2sb_io_in_r_valid; // @[NutShell.scala 62:16]
  assign io_frontend_r_bits_data = axi2sb_io_in_r_bits_data; // @[NutShell.scala 62:16]
  assign _T_4181 = nutcore__T_4181;
  assign _T_4184 = nutcore__T_4184;
  assign _T_4185 = nutcore__T_4185;
  assign falseWire = nutcore_falseWire;
  assign falseWire_0 = nutcore_falseWire_0;
  assign _T_4178 = nutcore__T_4178;
  assign _T_284_0 = nutcore__T_284_0;
  assign _T_284_1 = nutcore__T_284_1;
  assign _T_284_2 = nutcore__T_284_2;
  assign _T_284_3 = nutcore__T_284_3;
  assign _T_284_4 = nutcore__T_284_4;
  assign _T_284_5 = nutcore__T_284_5;
  assign _T_284_6 = nutcore__T_284_6;
  assign _T_284_7 = nutcore__T_284_7;
  assign _T_284_8 = nutcore__T_284_8;
  assign _T_284_9 = nutcore__T_284_9;
  assign _T_284_10 = nutcore__T_284_10;
  assign _T_284_11 = nutcore__T_284_11;
  assign _T_284_12 = nutcore__T_284_12;
  assign _T_284_13 = nutcore__T_284_13;
  assign _T_284_14 = nutcore__T_284_14;
  assign _T_284_15 = nutcore__T_284_15;
  assign _T_284_16 = nutcore__T_284_16;
  assign _T_284_17 = nutcore__T_284_17;
  assign _T_284_18 = nutcore__T_284_18;
  assign _T_284_19 = nutcore__T_284_19;
  assign _T_284_20 = nutcore__T_284_20;
  assign _T_284_21 = nutcore__T_284_21;
  assign _T_284_22 = nutcore__T_284_22;
  assign _T_284_23 = nutcore__T_284_23;
  assign _T_284_24 = nutcore__T_284_24;
  assign _T_284_25 = nutcore__T_284_25;
  assign _T_284_26 = nutcore__T_284_26;
  assign _T_284_27 = nutcore__T_284_27;
  assign _T_284_28 = nutcore__T_284_28;
  assign _T_284_29 = nutcore__T_284_29;
  assign _T_284_30 = nutcore__T_284_30;
  assign _T_284_31 = nutcore__T_284_31;
  assign _T_36 = nutcore__T_36_0;
  assign _T_32 = nutcore__T_32_0;
  assign _T_31 = nutcore__T_31_0;
  assign _T_37 = nutcore__T_37_0;
  assign _T_26 = nutcore__T_26_0;
  assign _T_4183 = nutcore__T_4183;
  assign _T_4182 = nutcore__T_4182;
  assign _T_33 = nutcore__T_33_0;
  assign _T_4179 = nutcore__T_4179;
  assign nutcore_clock = clock;
  assign nutcore_reset = reset;
  assign nutcore_io_imem_mem_req_ready = cohMg_io_in_req_ready; // @[NutShell.scala 56:15]
  assign nutcore_io_imem_mem_resp_valid = cohMg_io_in_resp_valid; // @[NutShell.scala 56:15]
  assign nutcore_io_imem_mem_resp_bits_cmd = cohMg_io_in_resp_bits_cmd; // @[NutShell.scala 56:15]
  assign nutcore_io_imem_mem_resp_bits_rdata = cohMg_io_in_resp_bits_rdata; // @[NutShell.scala 56:15]
  assign nutcore_io_dmem_mem_req_ready = xbar_io_in_1_req_ready; // @[NutShell.scala 59:17]
  assign nutcore_io_dmem_mem_resp_valid = xbar_io_in_1_resp_valid; // @[NutShell.scala 59:17]
  assign nutcore_io_dmem_mem_resp_bits_cmd = xbar_io_in_1_resp_bits_cmd; // @[NutShell.scala 59:17]
  assign nutcore_io_dmem_mem_resp_bits_rdata = xbar_io_in_1_resp_bits_rdata; // @[NutShell.scala 59:17]
  assign nutcore_io_dmem_coh_req_valid = cohMg_io_out_coh_req_valid; // @[NutShell.scala 57:23]
  assign nutcore_io_dmem_coh_req_bits_addr = cohMg_io_out_coh_req_bits_addr; // @[NutShell.scala 57:23]
  assign nutcore_io_dmem_coh_req_bits_wdata = cohMg_io_out_coh_req_bits_wdata; // @[NutShell.scala 57:23]
  assign nutcore_io_mmio_req_ready = mmioXbar_io_in_req_ready; // @[NutShell.scala 107:18]
  assign nutcore_io_mmio_resp_valid = mmioXbar_io_in_resp_valid; // @[NutShell.scala 107:18]
  assign nutcore_io_mmio_resp_bits_rdata = mmioXbar_io_in_resp_bits_rdata; // @[NutShell.scala 107:18]
  assign nutcore_io_frontend_req_valid = axi2sb_io_out_req_valid; // @[NutShell.scala 63:23]
  assign nutcore_io_frontend_req_bits_addr = axi2sb_io_out_req_bits_addr; // @[NutShell.scala 63:23]
  assign nutcore_io_frontend_req_bits_size = axi2sb_io_out_req_bits_size; // @[NutShell.scala 63:23]
  assign nutcore_io_frontend_req_bits_cmd = axi2sb_io_out_req_bits_cmd; // @[NutShell.scala 63:23]
  assign nutcore_io_frontend_req_bits_wmask = axi2sb_io_out_req_bits_wmask; // @[NutShell.scala 63:23]
  assign nutcore_io_frontend_req_bits_wdata = axi2sb_io_out_req_bits_wdata; // @[NutShell.scala 63:23]
  assign nutcore_io_frontend_resp_ready = axi2sb_io_out_resp_ready; // @[NutShell.scala 63:23]
  assign nutcore_io_extra_mtip = clint_io_extra_mtip;
  assign nutcore_DISPLAY_ENABLE = _T_13;
  assign nutcore_io_extra_meip_0 = plic_io_extra_meip_0;
  assign nutcore_io_extra_msip = clint_io_extra_msip;
  assign cohMg_clock = clock;
  assign cohMg_reset = reset;
  assign cohMg_io_in_req_valid = nutcore_io_imem_mem_req_valid; // @[NutShell.scala 56:15]
  assign cohMg_io_in_req_bits_addr = nutcore_io_imem_mem_req_bits_addr; // @[NutShell.scala 56:15]
  assign cohMg_io_in_req_bits_cmd = nutcore_io_imem_mem_req_bits_cmd; // @[NutShell.scala 56:15]
  assign cohMg_io_in_req_bits_wdata = nutcore_io_imem_mem_req_bits_wdata; // @[NutShell.scala 56:15]
  assign cohMg_io_out_mem_req_ready = xbar_io_in_0_req_ready; // @[NutShell.scala 58:17]
  assign cohMg_io_out_mem_resp_valid = xbar_io_in_0_resp_valid; // @[NutShell.scala 58:17]
  assign cohMg_io_out_mem_resp_bits_cmd = xbar_io_in_0_resp_bits_cmd; // @[NutShell.scala 58:17]
  assign cohMg_io_out_mem_resp_bits_rdata = xbar_io_in_0_resp_bits_rdata; // @[NutShell.scala 58:17]
  assign cohMg_io_out_coh_req_ready = nutcore_io_dmem_coh_req_ready; // @[NutShell.scala 57:23]
  assign cohMg_io_out_coh_resp_valid = nutcore_io_dmem_coh_resp_valid; // @[NutShell.scala 57:23]
  assign cohMg_io_out_coh_resp_bits_cmd = nutcore_io_dmem_coh_resp_bits_cmd; // @[NutShell.scala 57:23]
  assign cohMg_io_out_coh_resp_bits_rdata = nutcore_io_dmem_coh_resp_bits_rdata; // @[NutShell.scala 57:23]
  assign xbar_clock = clock;
  assign xbar_reset = reset;
  assign xbar_io_in_0_req_valid = cohMg_io_out_mem_req_valid; // @[NutShell.scala 58:17]
  assign xbar_io_in_0_req_bits_addr = cohMg_io_out_mem_req_bits_addr; // @[NutShell.scala 58:17]
  assign xbar_io_in_0_req_bits_cmd = cohMg_io_out_mem_req_bits_cmd; // @[NutShell.scala 58:17]
  assign xbar_io_in_0_req_bits_wmask = 8'hff; // @[NutShell.scala 58:17]
  assign xbar_io_in_0_req_bits_wdata = cohMg_io_out_mem_req_bits_wdata; // @[NutShell.scala 58:17]
  assign xbar_io_in_1_req_valid = nutcore_io_dmem_mem_req_valid; // @[NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_addr = nutcore_io_dmem_mem_req_bits_addr; // @[NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_size = 3'h3; // @[NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_cmd = nutcore_io_dmem_mem_req_bits_cmd; // @[NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_wmask = 8'hff; // @[NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_wdata = nutcore_io_dmem_mem_req_bits_wdata; // @[NutShell.scala 59:17]
  assign xbar_io_out_req_ready = Prefetcher_io_in_ready; // @[ToMemPort.scala 51:18 NutShell.scala 75:24]
  assign xbar_io_out_resp_valid = Cache_io_in_resp_valid; // @[ToMemPort.scala 51:18 NutShell.scala 77:24]
  assign xbar_io_out_resp_bits_cmd = Cache_io_in_resp_bits_cmd; // @[ToMemPort.scala 51:18 NutShell.scala 77:24]
  assign xbar_io_out_resp_bits_rdata = Cache_io_in_resp_bits_rdata; // @[ToMemPort.scala 51:18 NutShell.scala 77:24]
  assign axi2sb_clock = clock;
  assign axi2sb_reset = reset;
  assign axi2sb_io_in_aw_valid = io_frontend_aw_valid; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_aw_bits_addr = io_frontend_aw_bits_addr; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_aw_bits_len = io_frontend_aw_bits_len; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_aw_bits_size = io_frontend_aw_bits_size; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_w_valid = io_frontend_w_valid; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_w_bits_data = io_frontend_w_bits_data; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_w_bits_strb = io_frontend_w_bits_strb; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_b_ready = io_frontend_b_ready; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_ar_valid = io_frontend_ar_valid; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_ar_bits_addr = io_frontend_ar_bits_addr; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_r_ready = io_frontend_r_ready; // @[NutShell.scala 62:16]
  assign axi2sb_io_out_req_ready = nutcore_io_frontend_req_ready; // @[NutShell.scala 63:23]
  assign axi2sb_io_out_resp_valid = nutcore_io_frontend_resp_valid; // @[NutShell.scala 63:23]
  assign axi2sb_io_out_resp_bits_cmd = nutcore_io_frontend_resp_bits_cmd; // @[NutShell.scala 63:23]
  assign axi2sb_io_out_resp_bits_rdata = nutcore_io_frontend_resp_bits_rdata; // @[NutShell.scala 63:23]
  assign Prefetcher_clock = clock;
  assign Prefetcher_reset = reset;
  assign Prefetcher_io_in_valid = xbar_io_out_req_valid; // @[NutShell.scala 75:24]
  assign Prefetcher_io_in_bits_addr = xbar_io_out_req_bits_addr; // @[NutShell.scala 75:24]
  assign Prefetcher_io_in_bits_size = xbar_io_out_req_bits_size; // @[NutShell.scala 75:24]
  assign Prefetcher_io_in_bits_cmd = xbar_io_out_req_bits_cmd; // @[NutShell.scala 75:24]
  assign Prefetcher_io_in_bits_wmask = xbar_io_out_req_bits_wmask; // @[NutShell.scala 75:24]
  assign Prefetcher_io_in_bits_wdata = xbar_io_out_req_bits_wdata; // @[NutShell.scala 75:24]
  assign Prefetcher_io_out_ready = Cache_io_in_req_ready; // @[NutShell.scala 76:21]
  assign Prefetcher_DISPLAY_ENABLE = _T_13;
  assign Cache_clock = clock;
  assign Cache_reset = reset;
  assign Cache_io_in_req_valid = Prefetcher_io_out_valid; // @[Cache.scala 684:17]
  assign Cache_io_in_req_bits_addr = Prefetcher_io_out_bits_addr; // @[Cache.scala 684:17]
  assign Cache_io_in_req_bits_size = Prefetcher_io_out_bits_size; // @[Cache.scala 684:17]
  assign Cache_io_in_req_bits_cmd = Prefetcher_io_out_bits_cmd; // @[Cache.scala 684:17]
  assign Cache_io_in_req_bits_wmask = Prefetcher_io_out_bits_wmask; // @[Cache.scala 684:17]
  assign Cache_io_in_req_bits_wdata = Prefetcher_io_out_bits_wdata; // @[Cache.scala 684:17]
  assign Cache_io_out_mem_req_ready = memAddrMap_io_in_req_ready; // @[NutShell.scala 81:16]
  assign Cache_io_out_mem_resp_valid = memAddrMap_io_in_resp_valid; // @[NutShell.scala 81:16]
  assign Cache_io_out_mem_resp_bits_cmd = memAddrMap_io_in_resp_bits_cmd; // @[NutShell.scala 81:16]
  assign Cache_io_out_mem_resp_bits_rdata = memAddrMap_io_in_resp_bits_rdata; // @[NutShell.scala 81:16]
  assign Cache_DISPLAY_ENABLE = _T_13;
  assign memAddrMap_io_in_req_valid = Cache_io_out_mem_req_valid; // @[NutShell.scala 94:20]
  assign memAddrMap_io_in_req_bits_addr = Cache_io_out_mem_req_bits_addr; // @[NutShell.scala 94:20]
  assign memAddrMap_io_in_req_bits_cmd = Cache_io_out_mem_req_bits_cmd; // @[NutShell.scala 94:20]
  assign memAddrMap_io_in_req_bits_wdata = Cache_io_out_mem_req_bits_wdata; // @[NutShell.scala 94:20]
  assign memAddrMap_io_out_req_ready = SimpleBus2AXI4Converter_io_in_req_ready; // @[ToAXI4.scala 205:18]
  assign memAddrMap_io_out_resp_valid = SimpleBus2AXI4Converter_io_in_resp_valid; // @[ToAXI4.scala 205:18]
  assign memAddrMap_io_out_resp_bits_cmd = SimpleBus2AXI4Converter_io_in_resp_bits_cmd; // @[ToAXI4.scala 205:18]
  assign memAddrMap_io_out_resp_bits_rdata = SimpleBus2AXI4Converter_io_in_resp_bits_rdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_clock = clock;
  assign SimpleBus2AXI4Converter_reset = reset;
  assign SimpleBus2AXI4Converter_io_in_req_valid = memAddrMap_io_out_req_valid; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_io_in_req_bits_addr = memAddrMap_io_out_req_bits_addr; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_io_in_req_bits_cmd = memAddrMap_io_out_req_bits_cmd; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_io_in_req_bits_wdata = memAddrMap_io_out_req_bits_wdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_io_out_aw_ready = io_mem_aw_ready; // @[NutShell.scala 95:10]
  assign SimpleBus2AXI4Converter_io_out_w_ready = io_mem_w_ready; // @[NutShell.scala 95:10]
  assign SimpleBus2AXI4Converter_io_out_b_valid = io_mem_b_valid; // @[NutShell.scala 95:10]
  assign SimpleBus2AXI4Converter_io_out_ar_ready = io_mem_ar_ready; // @[NutShell.scala 95:10]
  assign SimpleBus2AXI4Converter_io_out_r_valid = io_mem_r_valid; // @[NutShell.scala 95:10]
  assign SimpleBus2AXI4Converter_io_out_r_bits_data = io_mem_r_bits_data; // @[NutShell.scala 95:10]
  assign SimpleBus2AXI4Converter_io_out_r_bits_last = io_mem_r_bits_last; // @[NutShell.scala 95:10]
  assign mmioXbar_clock = clock;
  assign mmioXbar_reset = reset;
  assign mmioXbar_io_in_req_valid = nutcore_io_mmio_req_valid; // @[NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_addr = nutcore_io_mmio_req_bits_addr; // @[NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_size = nutcore_io_mmio_req_bits_size; // @[NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_cmd = nutcore_io_mmio_req_bits_cmd; // @[NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_wmask = nutcore_io_mmio_req_bits_wmask; // @[NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_wdata = nutcore_io_mmio_req_bits_wdata; // @[NutShell.scala 107:18]
  assign mmioXbar_io_out_0_req_ready = io_mmio_req_ready; // @[NutShell.scala 111:18]
  assign mmioXbar_io_out_0_resp_valid = io_mmio_resp_valid; // @[NutShell.scala 111:18]
  assign mmioXbar_io_out_0_resp_bits_rdata = io_mmio_resp_bits_rdata; // @[NutShell.scala 111:18]
  assign mmioXbar_io_out_1_req_ready = SimpleBus2AXI4Converter_1_io_in_req_ready; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_1_resp_valid = SimpleBus2AXI4Converter_1_io_in_resp_valid; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_1_resp_bits_rdata = SimpleBus2AXI4Converter_1_io_in_resp_bits_rdata; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_2_req_ready = SimpleBus2AXI4Converter_2_io_in_req_ready; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_2_resp_valid = SimpleBus2AXI4Converter_2_io_in_resp_valid; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_2_resp_bits_rdata = SimpleBus2AXI4Converter_2_io_in_resp_bits_rdata; // @[ToAXI4.scala 205:18]
  assign mmioXbar_DISPLAY_ENABLE = _T_13;
  assign clint_clock = clock;
  assign clint_reset = reset;
  assign clint_io__in_aw_valid = SimpleBus2AXI4Converter_1_io_out_aw_valid; // @[NutShell.scala 114:15]
  assign clint_io__in_aw_bits_addr = SimpleBus2AXI4Converter_1_io_out_aw_bits_addr; // @[NutShell.scala 114:15]
  assign clint_io__in_w_valid = SimpleBus2AXI4Converter_1_io_out_w_valid; // @[NutShell.scala 114:15]
  assign clint_io__in_w_bits_data = SimpleBus2AXI4Converter_1_io_out_w_bits_data; // @[NutShell.scala 114:15]
  assign clint_io__in_w_bits_strb = SimpleBus2AXI4Converter_1_io_out_w_bits_strb; // @[NutShell.scala 114:15]
  assign clint_io__in_b_ready = SimpleBus2AXI4Converter_1_io_out_b_ready; // @[NutShell.scala 114:15]
  assign clint_io__in_ar_valid = SimpleBus2AXI4Converter_1_io_out_ar_valid; // @[NutShell.scala 114:15]
  assign clint_io__in_ar_bits_addr = SimpleBus2AXI4Converter_1_io_out_ar_bits_addr; // @[NutShell.scala 114:15]
  assign clint_io__in_r_ready = SimpleBus2AXI4Converter_1_io_out_r_ready; // @[NutShell.scala 114:15]
  assign clint_isWFI = nutcore__T_0;
  assign SimpleBus2AXI4Converter_1_clock = clock;
  assign SimpleBus2AXI4Converter_1_reset = reset;
  assign SimpleBus2AXI4Converter_1_io_in_req_valid = mmioXbar_io_out_1_req_valid; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_req_bits_addr = mmioXbar_io_out_1_req_bits_addr; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_req_bits_cmd = mmioXbar_io_out_1_req_bits_cmd; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_req_bits_wmask = mmioXbar_io_out_1_req_bits_wmask; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_req_bits_wdata = mmioXbar_io_out_1_req_bits_wdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_resp_ready = mmioXbar_io_out_1_resp_ready; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_out_aw_ready = clint_io__in_aw_ready; // @[NutShell.scala 114:15]
  assign SimpleBus2AXI4Converter_1_io_out_w_ready = clint_io__in_w_ready; // @[NutShell.scala 114:15]
  assign SimpleBus2AXI4Converter_1_io_out_b_valid = clint_io__in_b_valid; // @[NutShell.scala 114:15]
  assign SimpleBus2AXI4Converter_1_io_out_ar_ready = clint_io__in_ar_ready; // @[NutShell.scala 114:15]
  assign SimpleBus2AXI4Converter_1_io_out_r_valid = clint_io__in_r_valid; // @[NutShell.scala 114:15]
  assign SimpleBus2AXI4Converter_1_io_out_r_bits_data = clint_io__in_r_bits_data; // @[NutShell.scala 114:15]
  assign plic_clock = clock;
  assign plic_reset = reset;
  assign plic_io__in_aw_valid = SimpleBus2AXI4Converter_2_io_out_aw_valid; // @[NutShell.scala 121:14]
  assign plic_io__in_aw_bits_addr = SimpleBus2AXI4Converter_2_io_out_aw_bits_addr; // @[NutShell.scala 121:14]
  assign plic_io__in_w_valid = SimpleBus2AXI4Converter_2_io_out_w_valid; // @[NutShell.scala 121:14]
  assign plic_io__in_w_bits_data = SimpleBus2AXI4Converter_2_io_out_w_bits_data; // @[NutShell.scala 121:14]
  assign plic_io__in_w_bits_strb = SimpleBus2AXI4Converter_2_io_out_w_bits_strb; // @[NutShell.scala 121:14]
  assign plic_io__in_b_ready = SimpleBus2AXI4Converter_2_io_out_b_ready; // @[NutShell.scala 121:14]
  assign plic_io__in_ar_valid = SimpleBus2AXI4Converter_2_io_out_ar_valid; // @[NutShell.scala 121:14]
  assign plic_io__in_ar_bits_addr = SimpleBus2AXI4Converter_2_io_out_ar_bits_addr; // @[NutShell.scala 121:14]
  assign plic_io__in_r_ready = SimpleBus2AXI4Converter_2_io_out_r_ready; // @[NutShell.scala 121:14]
  assign plic_io__extra_intrVec = _T_5; // @[NutShell.scala 122:29]
  assign SimpleBus2AXI4Converter_2_clock = clock;
  assign SimpleBus2AXI4Converter_2_reset = reset;
  assign SimpleBus2AXI4Converter_2_io_in_req_valid = mmioXbar_io_out_2_req_valid; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_in_req_bits_addr = mmioXbar_io_out_2_req_bits_addr; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_in_req_bits_cmd = mmioXbar_io_out_2_req_bits_cmd; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_in_req_bits_wmask = mmioXbar_io_out_2_req_bits_wmask; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_in_req_bits_wdata = mmioXbar_io_out_2_req_bits_wdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_in_resp_ready = mmioXbar_io_out_2_resp_ready; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_out_aw_ready = plic_io__in_aw_ready; // @[NutShell.scala 121:14]
  assign SimpleBus2AXI4Converter_2_io_out_w_ready = plic_io__in_w_ready; // @[NutShell.scala 121:14]
  assign SimpleBus2AXI4Converter_2_io_out_b_valid = plic_io__in_b_valid; // @[NutShell.scala 121:14]
  assign SimpleBus2AXI4Converter_2_io_out_ar_ready = plic_io__in_ar_ready; // @[NutShell.scala 121:14]
  assign SimpleBus2AXI4Converter_2_io_out_r_valid = plic_io__in_r_valid; // @[NutShell.scala 121:14]
  assign SimpleBus2AXI4Converter_2_io_out_r_bits_data = plic_io__in_r_bits_data; // @[NutShell.scala 121:14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_4 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _T_5 = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_4 <= io_meip;
    _T_5 <= _T_4;
  end
endmodule
module AXI4RAM(
  input         clock,
  input         reset,
  output        io_in_aw_ready,
  input         io_in_aw_valid,
  input  [31:0] io_in_aw_bits_addr,
  output        io_in_w_ready,
  input         io_in_w_valid,
  input  [63:0] io_in_w_bits_data,
  input         io_in_w_bits_last,
  output        io_in_b_valid,
  output        io_in_ar_ready,
  input         io_in_ar_valid,
  input  [31:0] io_in_ar_bits_addr,
  input  [7:0]  io_in_ar_bits_len,
  input  [2:0]  io_in_ar_bits_size,
  input  [1:0]  io_in_ar_bits_burst,
  output        io_in_r_valid,
  output [63:0] io_in_r_bits_data,
  output        io_in_r_bits_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [63:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  RAMHelper_clk; // @[AXI4RAM.scala 52:21]
  wire [63:0] RAMHelper_rIdx; // @[AXI4RAM.scala 52:21]
  wire [63:0] RAMHelper_rdata; // @[AXI4RAM.scala 52:21]
  wire [63:0] RAMHelper_wIdx; // @[AXI4RAM.scala 52:21]
  wire [63:0] RAMHelper_wdata; // @[AXI4RAM.scala 52:21]
  wire [63:0] RAMHelper_wmask; // @[AXI4RAM.scala 52:21]
  wire  RAMHelper_wen; // @[AXI4RAM.scala 52:21]
  reg [7:0] value; // @[Counter.scala 29:33]
  reg [7:0] value_1; // @[Counter.scala 29:33]
  wire  _T_30 = io_in_ar_ready & io_in_ar_valid; // @[Decoupled.scala 40:37]
  reg [7:0] _T_32; // @[Reg.scala 27:20]
  wire [7:0] _GEN_0 = _T_30 ? io_in_ar_bits_len : _T_32; // @[Reg.scala 28:19]
  reg [1:0] _T_36; // @[Reg.scala 27:20]
  wire [1:0] _GEN_1 = _T_30 ? io_in_ar_bits_burst : _T_36; // @[Reg.scala 28:19]
  wire [31:0] _T_38 = {{24'd0}, io_in_ar_bits_len}; // @[AXI4Slave.scala 45:69 AXI4Slave.scala 45:69]
  wire [38:0] _GEN_24 = {{7'd0}, _T_38}; // @[AXI4Slave.scala 45:89]
  wire [38:0] _T_39 = _GEN_24 << io_in_ar_bits_size; // @[AXI4Slave.scala 45:89]
  wire [38:0] _T_40 = ~_T_39; // @[AXI4Slave.scala 45:42]
  wire [38:0] _GEN_25 = {{7'd0}, io_in_ar_bits_addr}; // @[AXI4Slave.scala 45:40]
  wire [38:0] _T_41 = _GEN_25 & _T_40; // @[AXI4Slave.scala 45:40]
  reg [38:0] _T_44; // @[Reg.scala 27:20]
  wire [38:0] _GEN_2 = _T_30 ? _T_41 : _T_44; // @[Reg.scala 28:19]
  wire [7:0] _T_49 = value_1 + 8'h1; // @[Counter.scala 39:22]
  wire  _T_50 = _GEN_1 == 2'h2; // @[AXI4Slave.scala 50:21]
  wire  _T_51 = value_1 == _GEN_0; // @[AXI4Slave.scala 50:68]
  wire  _T_52 = _T_50 & _T_51; // @[AXI4Slave.scala 50:51]
  wire [7:0] _GEN_3 = _T_52 ? 8'h0 : _T_49; // @[AXI4Slave.scala 50:77]
  reg  _T_79; // @[AXI4Slave.scala 73:17]
  wire  _T_81 = ~io_in_r_bits_last; // @[AXI4Slave.scala 73:65]
  wire  _T_82 = io_in_r_valid & _T_81; // @[AXI4Slave.scala 73:62]
  wire  ren = _T_79 | _T_82; // @[AXI4Slave.scala 73:46]
  wire [7:0] _GEN_4 = ren ? _GEN_3 : value_1; // @[AXI4Slave.scala 48:18]
  wire [7:0] _T_56 = value + 8'h1; // @[Counter.scala 39:22]
  wire [31:0] _T_58 = io_in_ar_bits_addr >> io_in_ar_bits_size; // @[AXI4Slave.scala 57:45]
  wire [31:0] _T_59 = _T_58 & _T_38; // @[AXI4Slave.scala 57:67]
  wire  _T_60 = io_in_ar_bits_len != 8'h0; // @[AXI4Slave.scala 58:32]
  wire  _T_61 = io_in_ar_bits_burst == 2'h2; // @[AXI4Slave.scala 58:62]
  wire  _T_62 = _T_60 & _T_61; // @[AXI4Slave.scala 58:40]
  wire  _T_63 = io_in_ar_bits_len == 8'h1; // @[AXI4Slave.scala 59:35]
  wire  _T_64 = io_in_ar_bits_len == 8'h3; // @[AXI4Slave.scala 59:63]
  wire  _T_65 = _T_63 | _T_64; // @[AXI4Slave.scala 59:43]
  wire  _T_66 = io_in_ar_bits_len == 8'h7; // @[AXI4Slave.scala 60:30]
  wire  _T_67 = _T_65 | _T_66; // @[AXI4Slave.scala 59:71]
  wire  _T_68 = io_in_ar_bits_len == 8'hf; // @[AXI4Slave.scala 60:58]
  wire  _T_69 = _T_67 | _T_68; // @[AXI4Slave.scala 60:38]
  wire  _T_71 = _T_69 | reset; // @[AXI4Slave.scala 59:17]
  wire  _T_72 = ~_T_71; // @[AXI4Slave.scala 59:17]
  wire [31:0] _GEN_7 = _T_30 ? _T_59 : {{24'd0}, _GEN_4}; // @[AXI4Slave.scala 56:29]
  wire  _T_75 = io_in_r_valid & io_in_r_bits_last; // @[AXI4Slave.scala 70:56]
  reg  r_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_8 = _T_75 ? 1'h0 : r_busy; // @[StopWatch.scala 26:19]
  wire  _GEN_9 = _T_30 | _GEN_8; // @[StopWatch.scala 27:20]
  wire  _T_85 = _T_30 | r_busy; // @[AXI4Slave.scala 74:52]
  wire  _T_86 = ren & _T_85; // @[AXI4Slave.scala 74:35]
  reg  _T_88; // @[StopWatch.scala 24:20]
  wire  _GEN_10 = io_in_r_valid ? 1'h0 : _T_88; // @[StopWatch.scala 26:19]
  wire  _GEN_11 = _T_86 | _GEN_10; // @[StopWatch.scala 27:20]
  reg [7:0] value_2; // @[Counter.scala 29:33]
  wire  _T_89 = io_in_aw_ready & io_in_aw_valid; // @[Decoupled.scala 40:37]
  reg [31:0] _T_91; // @[Reg.scala 27:20]
  wire [31:0] _GEN_12 = _T_89 ? io_in_aw_bits_addr : _T_91; // @[Reg.scala 28:19]
  wire  _T_93 = io_in_w_ready & io_in_w_valid; // @[Decoupled.scala 40:37]
  wire [7:0] _T_96 = value_2 + 8'h1; // @[Counter.scala 39:22]
  reg  w_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_15 = io_in_b_valid ? 1'h0 : w_busy; // @[StopWatch.scala 26:19]
  wire  _GEN_16 = _T_89 | _GEN_15; // @[StopWatch.scala 27:20]
  wire  _T_102 = _T_93 & io_in_w_bits_last; // @[AXI4Slave.scala 97:43]
  reg  _T_104; // @[StopWatch.scala 24:20]
  wire  _GEN_17 = io_in_b_valid ? 1'h0 : _T_104; // @[StopWatch.scala 26:19]
  wire  _GEN_18 = _T_102 | _GEN_17; // @[StopWatch.scala 27:20]
  wire [31:0] _T_113 = _GEN_12 & 32'h7ffffff; // @[AXI4RAM.scala 44:33]
  wire [28:0] _GEN_27 = {{21'd0}, value_2}; // @[AXI4RAM.scala 47:27]
  wire [28:0] wIdx = _T_113[31:3] + _GEN_27; // @[AXI4RAM.scala 47:27]
  wire [38:0] _T_116 = _GEN_2 & 39'h7ffffff; // @[AXI4RAM.scala 44:33]
  wire [35:0] _GEN_28 = {{28'd0}, value_1}; // @[AXI4RAM.scala 48:27]
  wire [35:0] rIdx = _T_116[38:3] + _GEN_28; // @[AXI4RAM.scala 48:27]
  wire  _T_120 = wIdx < 29'h1000000; // @[AXI4RAM.scala 45:32]
  reg [63:0] _T_121; // @[Reg.scala 15:16]
  wire  _GEN_31 = _T_30 & _T_62; // @[AXI4Slave.scala 59:17]
  RAMHelper RAMHelper ( // @[AXI4RAM.scala 52:21]
    .clk(RAMHelper_clk),
    .rIdx(RAMHelper_rIdx),
    .rdata(RAMHelper_rdata),
    .wIdx(RAMHelper_wIdx),
    .wdata(RAMHelper_wdata),
    .wmask(RAMHelper_wmask),
    .wen(RAMHelper_wen)
  );
  assign io_in_aw_ready = ~w_busy; // @[AXI4Slave.scala 94:15]
  assign io_in_w_ready = io_in_aw_valid | w_busy; // @[AXI4Slave.scala 95:15]
  assign io_in_b_valid = _T_104; // @[AXI4Slave.scala 97:14]
  assign io_in_ar_ready = 1'h1; // @[AXI4Slave.scala 71:15]
  assign io_in_r_valid = _T_88; // @[AXI4Slave.scala 74:14]
  assign io_in_r_bits_data = _T_121; // @[AXI4RAM.scala 69:18]
  assign io_in_r_bits_last = value == _GEN_0; // @[AXI4Slave.scala 47:24]
  assign RAMHelper_clk = clock; // @[AXI4RAM.scala 53:16]
  assign RAMHelper_rIdx = {{28'd0}, rIdx}; // @[AXI4RAM.scala 54:17]
  assign RAMHelper_wIdx = {{35'd0}, wIdx}; // @[AXI4RAM.scala 55:17]
  assign RAMHelper_wdata = io_in_w_bits_data; // @[AXI4RAM.scala 56:18]
  assign RAMHelper_wmask = 64'hffffffffffffffff; // @[AXI4RAM.scala 57:18]
  assign RAMHelper_wen = _T_93 & _T_120; // @[AXI4RAM.scala 58:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  value_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  _T_32 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  _T_36 = _RAND_3[1:0];
  _RAND_4 = {2{`RANDOM}};
  _T_44 = _RAND_4[38:0];
  _RAND_5 = {1{`RANDOM}};
  _T_79 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  r_busy = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_88 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  value_2 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  _T_91 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  w_busy = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _T_104 = _RAND_11[0:0];
  _RAND_12 = {2{`RANDOM}};
  _T_121 = _RAND_12[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 8'h0;
    end else if (io_in_r_valid) begin
      if (io_in_r_bits_last) begin
        value <= 8'h0;
      end else begin
        value <= _T_56;
      end
    end
    if (reset) begin
      value_1 <= 8'h0;
    end else begin
      value_1 <= _GEN_7[7:0];
    end
    if (reset) begin
      _T_32 <= 8'h0;
    end else if (_T_30) begin
      _T_32 <= io_in_ar_bits_len;
    end
    if (reset) begin
      _T_36 <= 2'h0;
    end else if (_T_30) begin
      _T_36 <= io_in_ar_bits_burst;
    end
    if (reset) begin
      _T_44 <= 39'h0;
    end else if (_T_30) begin
      _T_44 <= _T_41;
    end
    if (reset) begin
      _T_79 <= 1'h0;
    end else begin
      _T_79 <= _T_30;
    end
    if (reset) begin
      r_busy <= 1'h0;
    end else begin
      r_busy <= _GEN_9;
    end
    if (reset) begin
      _T_88 <= 1'h0;
    end else begin
      _T_88 <= _GEN_11;
    end
    if (reset) begin
      value_2 <= 8'h0;
    end else if (_T_93) begin
      if (io_in_w_bits_last) begin
        value_2 <= 8'h0;
      end else begin
        value_2 <= _T_96;
      end
    end
    if (reset) begin
      _T_91 <= 32'h0;
    end else if (_T_89) begin
      _T_91 <= io_in_aw_bits_addr;
    end
    if (reset) begin
      w_busy <= 1'h0;
    end else begin
      w_busy <= _GEN_16;
    end
    if (reset) begin
      _T_104 <= 1'h0;
    end else begin
      _T_104 <= _GEN_18;
    end
    if (ren) begin
      _T_121 <= RAMHelper_rdata;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_31 & _T_72) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4Slave.scala:59 assert(axi4.ar.bits.len === 1.U || axi4.ar.bits.len === 3.U ||\n"); // @[AXI4Slave.scala 59:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_31 & _T_72) begin
          $fatal; // @[AXI4Slave.scala 59:17]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module LatencyPipe(
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [7:0]  io_in_bits_len,
  input  [2:0]  io_in_bits_size,
  input  [1:0]  io_in_bits_burst,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [7:0]  io_out_bits_len,
  output [2:0]  io_out_bits_size,
  output [1:0]  io_out_bits_burst
);
  assign io_in_ready = io_out_ready; // @[LatencyPipe.scala 16:10]
  assign io_out_valid = io_in_valid; // @[LatencyPipe.scala 16:10]
  assign io_out_bits_addr = io_in_bits_addr; // @[LatencyPipe.scala 16:10]
  assign io_out_bits_len = io_in_bits_len; // @[LatencyPipe.scala 16:10]
  assign io_out_bits_size = io_in_bits_size; // @[LatencyPipe.scala 16:10]
  assign io_out_bits_burst = io_in_bits_burst; // @[LatencyPipe.scala 16:10]
endmodule
module AXI4Delayer(
  output        io_in_aw_ready,
  input         io_in_aw_valid,
  input  [31:0] io_in_aw_bits_addr,
  input  [7:0]  io_in_aw_bits_len,
  input  [2:0]  io_in_aw_bits_size,
  input  [1:0]  io_in_aw_bits_burst,
  output        io_in_w_ready,
  input         io_in_w_valid,
  input  [63:0] io_in_w_bits_data,
  input         io_in_w_bits_last,
  output        io_in_b_valid,
  output        io_in_ar_ready,
  input         io_in_ar_valid,
  input  [31:0] io_in_ar_bits_addr,
  input  [7:0]  io_in_ar_bits_len,
  output        io_in_r_valid,
  output [63:0] io_in_r_bits_data,
  output        io_in_r_bits_last,
  input         io_out_aw_ready,
  output        io_out_aw_valid,
  output [31:0] io_out_aw_bits_addr,
  input         io_out_w_ready,
  output        io_out_w_valid,
  output [63:0] io_out_w_bits_data,
  output        io_out_w_bits_last,
  input         io_out_b_valid,
  output        io_out_ar_valid,
  output [31:0] io_out_ar_bits_addr,
  output [7:0]  io_out_ar_bits_len,
  output [2:0]  io_out_ar_bits_size,
  output [1:0]  io_out_ar_bits_burst,
  input         io_out_r_valid,
  input  [63:0] io_out_r_bits_data,
  input         io_out_r_bits_last
);
  wire  LatencyPipe_io_in_ready; // @[LatencyPipe.scala 21:22]
  wire  LatencyPipe_io_in_valid; // @[LatencyPipe.scala 21:22]
  wire [31:0] LatencyPipe_io_in_bits_addr; // @[LatencyPipe.scala 21:22]
  wire [7:0] LatencyPipe_io_in_bits_len; // @[LatencyPipe.scala 21:22]
  wire [2:0] LatencyPipe_io_in_bits_size; // @[LatencyPipe.scala 21:22]
  wire [1:0] LatencyPipe_io_in_bits_burst; // @[LatencyPipe.scala 21:22]
  wire  LatencyPipe_io_out_ready; // @[LatencyPipe.scala 21:22]
  wire  LatencyPipe_io_out_valid; // @[LatencyPipe.scala 21:22]
  wire [31:0] LatencyPipe_io_out_bits_addr; // @[LatencyPipe.scala 21:22]
  wire [7:0] LatencyPipe_io_out_bits_len; // @[LatencyPipe.scala 21:22]
  wire [2:0] LatencyPipe_io_out_bits_size; // @[LatencyPipe.scala 21:22]
  wire [1:0] LatencyPipe_io_out_bits_burst; // @[LatencyPipe.scala 21:22]
  wire  LatencyPipe_1_io_in_ready; // @[LatencyPipe.scala 21:22]
  wire  LatencyPipe_1_io_in_valid; // @[LatencyPipe.scala 21:22]
  wire [31:0] LatencyPipe_1_io_in_bits_addr; // @[LatencyPipe.scala 21:22]
  wire [7:0] LatencyPipe_1_io_in_bits_len; // @[LatencyPipe.scala 21:22]
  wire [2:0] LatencyPipe_1_io_in_bits_size; // @[LatencyPipe.scala 21:22]
  wire [1:0] LatencyPipe_1_io_in_bits_burst; // @[LatencyPipe.scala 21:22]
  wire  LatencyPipe_1_io_out_ready; // @[LatencyPipe.scala 21:22]
  wire  LatencyPipe_1_io_out_valid; // @[LatencyPipe.scala 21:22]
  wire [31:0] LatencyPipe_1_io_out_bits_addr; // @[LatencyPipe.scala 21:22]
  wire [7:0] LatencyPipe_1_io_out_bits_len; // @[LatencyPipe.scala 21:22]
  wire [2:0] LatencyPipe_1_io_out_bits_size; // @[LatencyPipe.scala 21:22]
  wire [1:0] LatencyPipe_1_io_out_bits_burst; // @[LatencyPipe.scala 21:22]
  LatencyPipe LatencyPipe ( // @[LatencyPipe.scala 21:22]
    .io_in_ready(LatencyPipe_io_in_ready),
    .io_in_valid(LatencyPipe_io_in_valid),
    .io_in_bits_addr(LatencyPipe_io_in_bits_addr),
    .io_in_bits_len(LatencyPipe_io_in_bits_len),
    .io_in_bits_size(LatencyPipe_io_in_bits_size),
    .io_in_bits_burst(LatencyPipe_io_in_bits_burst),
    .io_out_ready(LatencyPipe_io_out_ready),
    .io_out_valid(LatencyPipe_io_out_valid),
    .io_out_bits_addr(LatencyPipe_io_out_bits_addr),
    .io_out_bits_len(LatencyPipe_io_out_bits_len),
    .io_out_bits_size(LatencyPipe_io_out_bits_size),
    .io_out_bits_burst(LatencyPipe_io_out_bits_burst)
  );
  LatencyPipe LatencyPipe_1 ( // @[LatencyPipe.scala 21:22]
    .io_in_ready(LatencyPipe_1_io_in_ready),
    .io_in_valid(LatencyPipe_1_io_in_valid),
    .io_in_bits_addr(LatencyPipe_1_io_in_bits_addr),
    .io_in_bits_len(LatencyPipe_1_io_in_bits_len),
    .io_in_bits_size(LatencyPipe_1_io_in_bits_size),
    .io_in_bits_burst(LatencyPipe_1_io_in_bits_burst),
    .io_out_ready(LatencyPipe_1_io_out_ready),
    .io_out_valid(LatencyPipe_1_io_out_valid),
    .io_out_bits_addr(LatencyPipe_1_io_out_bits_addr),
    .io_out_bits_len(LatencyPipe_1_io_out_bits_len),
    .io_out_bits_size(LatencyPipe_1_io_out_bits_size),
    .io_out_bits_burst(LatencyPipe_1_io_out_bits_burst)
  );
  assign io_in_aw_ready = LatencyPipe_1_io_in_ready; // @[LatencyPipe.scala 22:16]
  assign io_in_w_ready = io_out_w_ready; // @[Delayer.scala 17:13]
  assign io_in_b_valid = io_out_b_valid; // @[Delayer.scala 18:13]
  assign io_in_ar_ready = LatencyPipe_io_in_ready; // @[LatencyPipe.scala 22:16]
  assign io_in_r_valid = io_out_r_valid; // @[Delayer.scala 19:13]
  assign io_in_r_bits_data = io_out_r_bits_data; // @[Delayer.scala 19:13]
  assign io_in_r_bits_last = io_out_r_bits_last; // @[Delayer.scala 19:13]
  assign io_out_aw_valid = LatencyPipe_1_io_out_valid; // @[Delayer.scala 16:13]
  assign io_out_aw_bits_addr = LatencyPipe_1_io_out_bits_addr; // @[Delayer.scala 16:13]
  assign io_out_w_valid = io_in_w_valid; // @[Delayer.scala 17:13]
  assign io_out_w_bits_data = io_in_w_bits_data; // @[Delayer.scala 17:13]
  assign io_out_w_bits_last = io_in_w_bits_last; // @[Delayer.scala 17:13]
  assign io_out_ar_valid = LatencyPipe_io_out_valid; // @[Delayer.scala 15:13]
  assign io_out_ar_bits_addr = LatencyPipe_io_out_bits_addr; // @[Delayer.scala 15:13]
  assign io_out_ar_bits_len = LatencyPipe_io_out_bits_len; // @[Delayer.scala 15:13]
  assign io_out_ar_bits_size = LatencyPipe_io_out_bits_size; // @[Delayer.scala 15:13]
  assign io_out_ar_bits_burst = LatencyPipe_io_out_bits_burst; // @[Delayer.scala 15:13]
  assign LatencyPipe_io_in_valid = io_in_ar_valid; // @[LatencyPipe.scala 22:16]
  assign LatencyPipe_io_in_bits_addr = io_in_ar_bits_addr; // @[LatencyPipe.scala 22:16]
  assign LatencyPipe_io_in_bits_len = io_in_ar_bits_len; // @[LatencyPipe.scala 22:16]
  assign LatencyPipe_io_in_bits_size = 3'h3; // @[LatencyPipe.scala 22:16]
  assign LatencyPipe_io_in_bits_burst = 2'h2; // @[LatencyPipe.scala 22:16]
  assign LatencyPipe_io_out_ready = 1'h1; // @[Delayer.scala 15:13]
  assign LatencyPipe_1_io_in_valid = io_in_aw_valid; // @[LatencyPipe.scala 22:16]
  assign LatencyPipe_1_io_in_bits_addr = io_in_aw_bits_addr; // @[LatencyPipe.scala 22:16]
  assign LatencyPipe_1_io_in_bits_len = io_in_aw_bits_len; // @[LatencyPipe.scala 22:16]
  assign LatencyPipe_1_io_in_bits_size = io_in_aw_bits_size; // @[LatencyPipe.scala 22:16]
  assign LatencyPipe_1_io_in_bits_burst = io_in_aw_bits_burst; // @[LatencyPipe.scala 22:16]
  assign LatencyPipe_1_io_out_ready = io_out_aw_ready; // @[Delayer.scala 16:13]
endmodule
module SimpleBusCrossbar1toN_1(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [2:0]  io_in_req_bits_size,
  input  [3:0]  io_in_req_bits_cmd,
  input  [7:0]  io_in_req_bits_wmask,
  input  [63:0] io_in_req_bits_wdata,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_0_req_ready,
  output        io_out_0_req_valid,
  output [31:0] io_out_0_req_bits_addr,
  output [2:0]  io_out_0_req_bits_size,
  output [3:0]  io_out_0_req_bits_cmd,
  output [7:0]  io_out_0_req_bits_wmask,
  output [63:0] io_out_0_req_bits_wdata,
  output        io_out_0_resp_ready,
  input         io_out_0_resp_valid,
  input  [63:0] io_out_0_resp_bits_rdata,
  input         io_out_1_req_ready,
  output        io_out_1_req_valid,
  output [31:0] io_out_1_req_bits_addr,
  output [2:0]  io_out_1_req_bits_size,
  output [3:0]  io_out_1_req_bits_cmd,
  output [7:0]  io_out_1_req_bits_wmask,
  output [63:0] io_out_1_req_bits_wdata,
  output        io_out_1_resp_ready,
  input         io_out_1_resp_valid,
  input  [63:0] io_out_1_resp_bits_rdata,
  input         io_out_2_req_ready,
  output        io_out_2_req_valid,
  output [31:0] io_out_2_req_bits_addr,
  output [2:0]  io_out_2_req_bits_size,
  output [3:0]  io_out_2_req_bits_cmd,
  output [7:0]  io_out_2_req_bits_wmask,
  output [63:0] io_out_2_req_bits_wdata,
  output        io_out_2_resp_ready,
  input         io_out_2_resp_valid,
  input  [63:0] io_out_2_resp_bits_rdata,
  input         io_out_3_req_ready,
  output        io_out_3_req_valid,
  output [31:0] io_out_3_req_bits_addr,
  output [2:0]  io_out_3_req_bits_size,
  output [3:0]  io_out_3_req_bits_cmd,
  output [7:0]  io_out_3_req_bits_wmask,
  output [63:0] io_out_3_req_bits_wdata,
  output        io_out_3_resp_ready,
  input         io_out_3_resp_valid,
  input  [63:0] io_out_3_resp_bits_rdata,
  input         io_out_4_req_ready,
  output        io_out_4_req_valid,
  output [31:0] io_out_4_req_bits_addr,
  output [2:0]  io_out_4_req_bits_size,
  output [3:0]  io_out_4_req_bits_cmd,
  output [7:0]  io_out_4_req_bits_wmask,
  output [63:0] io_out_4_req_bits_wdata,
  output        io_out_4_resp_ready,
  input         io_out_4_resp_valid,
  input  [63:0] io_out_4_resp_bits_rdata,
  input         io_out_5_req_ready,
  output        io_out_5_req_valid,
  output [31:0] io_out_5_req_bits_addr,
  output [2:0]  io_out_5_req_bits_size,
  output [3:0]  io_out_5_req_bits_cmd,
  output [7:0]  io_out_5_req_bits_wmask,
  output [63:0] io_out_5_req_bits_wdata,
  output        io_out_5_resp_ready,
  input         io_out_5_resp_valid,
  input  [63:0] io_out_5_resp_bits_rdata,
  input         io_out_6_req_ready,
  output        io_out_6_req_valid,
  output [31:0] io_out_6_req_bits_addr,
  output [2:0]  io_out_6_req_bits_size,
  output [3:0]  io_out_6_req_bits_cmd,
  output [7:0]  io_out_6_req_bits_wmask,
  output [63:0] io_out_6_req_bits_wdata,
  output        io_out_6_resp_ready,
  input         io_out_6_resp_valid,
  input  [63:0] io_out_6_resp_bits_rdata,
  input         io_out_7_req_ready,
  output        io_out_7_req_valid,
  output [31:0] io_out_7_req_bits_addr,
  output [2:0]  io_out_7_req_bits_size,
  output [3:0]  io_out_7_req_bits_cmd,
  output [7:0]  io_out_7_req_bits_wmask,
  output [63:0] io_out_7_req_bits_wdata,
  output        io_out_7_resp_ready,
  input         io_out_7_resp_valid,
  input  [63:0] io_out_7_resp_bits_rdata,
  input         DISPLAY_ENABLE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[Crossbar.scala 31:22]
  wire  _T = io_in_req_bits_addr >= 32'h40600000; // @[Crossbar.scala 36:20]
  wire  _T_1 = io_in_req_bits_addr < 32'h40600010; // @[Crossbar.scala 36:42]
  wire  outSelVec_0 = _T & _T_1; // @[Crossbar.scala 36:34]
  wire  _T_3 = io_in_req_bits_addr >= 32'h50000000; // @[Crossbar.scala 36:20]
  wire  _T_4 = io_in_req_bits_addr < 32'h50400000; // @[Crossbar.scala 36:42]
  wire  outSelVec_1 = _T_3 & _T_4; // @[Crossbar.scala 36:34]
  wire  _T_6 = io_in_req_bits_addr >= 32'h40001000; // @[Crossbar.scala 36:20]
  wire  _T_7 = io_in_req_bits_addr < 32'h40001008; // @[Crossbar.scala 36:42]
  wire  outSelVec_2 = _T_6 & _T_7; // @[Crossbar.scala 36:34]
  wire  _T_9 = io_in_req_bits_addr >= 32'h40000000; // @[Crossbar.scala 36:20]
  wire  _T_10 = io_in_req_bits_addr < 32'h40001000; // @[Crossbar.scala 36:42]
  wire  outSelVec_3 = _T_9 & _T_10; // @[Crossbar.scala 36:34]
  wire  _T_12 = io_in_req_bits_addr >= 32'h40002000; // @[Crossbar.scala 36:20]
  wire  _T_13 = io_in_req_bits_addr < 32'h40003000; // @[Crossbar.scala 36:42]
  wire  outSelVec_4 = _T_12 & _T_13; // @[Crossbar.scala 36:34]
  wire  _T_15 = io_in_req_bits_addr >= 32'h42000000; // @[Crossbar.scala 36:20]
  wire  _T_16 = io_in_req_bits_addr < 32'h42001000; // @[Crossbar.scala 36:42]
  wire  outSelVec_5 = _T_15 & _T_16; // @[Crossbar.scala 36:34]
  wire  _T_18 = io_in_req_bits_addr >= 32'h40004000; // @[Crossbar.scala 36:20]
  wire  _T_19 = io_in_req_bits_addr < 32'h40005000; // @[Crossbar.scala 36:42]
  wire  outSelVec_6 = _T_18 & _T_19; // @[Crossbar.scala 36:34]
  wire  _T_21 = io_in_req_bits_addr >= 32'h40003000; // @[Crossbar.scala 36:20]
  wire  _T_22 = io_in_req_bits_addr < 32'h40004000; // @[Crossbar.scala 36:42]
  wire  outSelVec_7 = _T_21 & _T_22; // @[Crossbar.scala 36:34]
  wire [2:0] _T_24 = outSelVec_6 ? 3'h6 : 3'h7; // @[Mux.scala 47:69]
  wire [2:0] _T_25 = outSelVec_5 ? 3'h5 : _T_24; // @[Mux.scala 47:69]
  wire [2:0] _T_26 = outSelVec_4 ? 3'h4 : _T_25; // @[Mux.scala 47:69]
  wire [2:0] _T_27 = outSelVec_3 ? 3'h3 : _T_26; // @[Mux.scala 47:69]
  wire [2:0] _T_28 = outSelVec_2 ? 3'h2 : _T_27; // @[Mux.scala 47:69]
  wire [2:0] _T_29 = outSelVec_1 ? 3'h1 : _T_28; // @[Mux.scala 47:69]
  wire [2:0] outSelIdx = outSelVec_0 ? 3'h0 : _T_29; // @[Mux.scala 47:69]
  wire  _GEN_11 = 3'h1 == outSelIdx ? io_out_1_req_ready : io_out_0_req_ready; // @[Decoupled.scala 40:37]
  wire  _GEN_12 = 3'h1 == outSelIdx ? io_out_1_req_valid : io_out_0_req_valid; // @[Decoupled.scala 40:37]
  wire [31:0] _GEN_13 = 3'h1 == outSelIdx ? io_out_1_req_bits_addr : io_out_0_req_bits_addr; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_14 = 3'h1 == outSelIdx ? io_out_1_req_bits_size : io_out_0_req_bits_size; // @[Decoupled.scala 40:37]
  wire [3:0] _GEN_15 = 3'h1 == outSelIdx ? io_out_1_req_bits_cmd : io_out_0_req_bits_cmd; // @[Decoupled.scala 40:37]
  wire [7:0] _GEN_16 = 3'h1 == outSelIdx ? io_out_1_req_bits_wmask : io_out_0_req_bits_wmask; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_17 = 3'h1 == outSelIdx ? io_out_1_req_bits_wdata : io_out_0_req_bits_wdata; // @[Decoupled.scala 40:37]
  wire  _GEN_18 = 3'h1 == outSelIdx ? io_out_1_resp_ready : io_out_0_resp_ready; // @[Decoupled.scala 40:37]
  wire  _GEN_19 = 3'h1 == outSelIdx ? io_out_1_resp_valid : io_out_0_resp_valid; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_21 = 3'h1 == outSelIdx ? io_out_1_resp_bits_rdata : io_out_0_resp_bits_rdata; // @[Decoupled.scala 40:37]
  wire  _GEN_22 = 3'h2 == outSelIdx ? io_out_2_req_ready : _GEN_11; // @[Decoupled.scala 40:37]
  wire  _GEN_23 = 3'h2 == outSelIdx ? io_out_2_req_valid : _GEN_12; // @[Decoupled.scala 40:37]
  wire [31:0] _GEN_24 = 3'h2 == outSelIdx ? io_out_2_req_bits_addr : _GEN_13; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_25 = 3'h2 == outSelIdx ? io_out_2_req_bits_size : _GEN_14; // @[Decoupled.scala 40:37]
  wire [3:0] _GEN_26 = 3'h2 == outSelIdx ? io_out_2_req_bits_cmd : _GEN_15; // @[Decoupled.scala 40:37]
  wire [7:0] _GEN_27 = 3'h2 == outSelIdx ? io_out_2_req_bits_wmask : _GEN_16; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_28 = 3'h2 == outSelIdx ? io_out_2_req_bits_wdata : _GEN_17; // @[Decoupled.scala 40:37]
  wire  _GEN_29 = 3'h2 == outSelIdx ? io_out_2_resp_ready : _GEN_18; // @[Decoupled.scala 40:37]
  wire  _GEN_30 = 3'h2 == outSelIdx ? io_out_2_resp_valid : _GEN_19; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_32 = 3'h2 == outSelIdx ? io_out_2_resp_bits_rdata : _GEN_21; // @[Decoupled.scala 40:37]
  wire  _GEN_33 = 3'h3 == outSelIdx ? io_out_3_req_ready : _GEN_22; // @[Decoupled.scala 40:37]
  wire  _GEN_34 = 3'h3 == outSelIdx ? io_out_3_req_valid : _GEN_23; // @[Decoupled.scala 40:37]
  wire [31:0] _GEN_35 = 3'h3 == outSelIdx ? io_out_3_req_bits_addr : _GEN_24; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_36 = 3'h3 == outSelIdx ? io_out_3_req_bits_size : _GEN_25; // @[Decoupled.scala 40:37]
  wire [3:0] _GEN_37 = 3'h3 == outSelIdx ? io_out_3_req_bits_cmd : _GEN_26; // @[Decoupled.scala 40:37]
  wire [7:0] _GEN_38 = 3'h3 == outSelIdx ? io_out_3_req_bits_wmask : _GEN_27; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_39 = 3'h3 == outSelIdx ? io_out_3_req_bits_wdata : _GEN_28; // @[Decoupled.scala 40:37]
  wire  _GEN_40 = 3'h3 == outSelIdx ? io_out_3_resp_ready : _GEN_29; // @[Decoupled.scala 40:37]
  wire  _GEN_41 = 3'h3 == outSelIdx ? io_out_3_resp_valid : _GEN_30; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_43 = 3'h3 == outSelIdx ? io_out_3_resp_bits_rdata : _GEN_32; // @[Decoupled.scala 40:37]
  wire  _GEN_44 = 3'h4 == outSelIdx ? io_out_4_req_ready : _GEN_33; // @[Decoupled.scala 40:37]
  wire  _GEN_45 = 3'h4 == outSelIdx ? io_out_4_req_valid : _GEN_34; // @[Decoupled.scala 40:37]
  wire [31:0] _GEN_46 = 3'h4 == outSelIdx ? io_out_4_req_bits_addr : _GEN_35; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_47 = 3'h4 == outSelIdx ? io_out_4_req_bits_size : _GEN_36; // @[Decoupled.scala 40:37]
  wire [3:0] _GEN_48 = 3'h4 == outSelIdx ? io_out_4_req_bits_cmd : _GEN_37; // @[Decoupled.scala 40:37]
  wire [7:0] _GEN_49 = 3'h4 == outSelIdx ? io_out_4_req_bits_wmask : _GEN_38; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_50 = 3'h4 == outSelIdx ? io_out_4_req_bits_wdata : _GEN_39; // @[Decoupled.scala 40:37]
  wire  _GEN_51 = 3'h4 == outSelIdx ? io_out_4_resp_ready : _GEN_40; // @[Decoupled.scala 40:37]
  wire  _GEN_52 = 3'h4 == outSelIdx ? io_out_4_resp_valid : _GEN_41; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_54 = 3'h4 == outSelIdx ? io_out_4_resp_bits_rdata : _GEN_43; // @[Decoupled.scala 40:37]
  wire  _GEN_55 = 3'h5 == outSelIdx ? io_out_5_req_ready : _GEN_44; // @[Decoupled.scala 40:37]
  wire  _GEN_56 = 3'h5 == outSelIdx ? io_out_5_req_valid : _GEN_45; // @[Decoupled.scala 40:37]
  wire [31:0] _GEN_57 = 3'h5 == outSelIdx ? io_out_5_req_bits_addr : _GEN_46; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_58 = 3'h5 == outSelIdx ? io_out_5_req_bits_size : _GEN_47; // @[Decoupled.scala 40:37]
  wire [3:0] _GEN_59 = 3'h5 == outSelIdx ? io_out_5_req_bits_cmd : _GEN_48; // @[Decoupled.scala 40:37]
  wire [7:0] _GEN_60 = 3'h5 == outSelIdx ? io_out_5_req_bits_wmask : _GEN_49; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_61 = 3'h5 == outSelIdx ? io_out_5_req_bits_wdata : _GEN_50; // @[Decoupled.scala 40:37]
  wire  _GEN_62 = 3'h5 == outSelIdx ? io_out_5_resp_ready : _GEN_51; // @[Decoupled.scala 40:37]
  wire  _GEN_63 = 3'h5 == outSelIdx ? io_out_5_resp_valid : _GEN_52; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_65 = 3'h5 == outSelIdx ? io_out_5_resp_bits_rdata : _GEN_54; // @[Decoupled.scala 40:37]
  wire  _GEN_66 = 3'h6 == outSelIdx ? io_out_6_req_ready : _GEN_55; // @[Decoupled.scala 40:37]
  wire  _GEN_67 = 3'h6 == outSelIdx ? io_out_6_req_valid : _GEN_56; // @[Decoupled.scala 40:37]
  wire [31:0] _GEN_68 = 3'h6 == outSelIdx ? io_out_6_req_bits_addr : _GEN_57; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_69 = 3'h6 == outSelIdx ? io_out_6_req_bits_size : _GEN_58; // @[Decoupled.scala 40:37]
  wire [3:0] _GEN_70 = 3'h6 == outSelIdx ? io_out_6_req_bits_cmd : _GEN_59; // @[Decoupled.scala 40:37]
  wire [7:0] _GEN_71 = 3'h6 == outSelIdx ? io_out_6_req_bits_wmask : _GEN_60; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_72 = 3'h6 == outSelIdx ? io_out_6_req_bits_wdata : _GEN_61; // @[Decoupled.scala 40:37]
  wire  _GEN_73 = 3'h6 == outSelIdx ? io_out_6_resp_ready : _GEN_62; // @[Decoupled.scala 40:37]
  wire  _GEN_74 = 3'h6 == outSelIdx ? io_out_6_resp_valid : _GEN_63; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_76 = 3'h6 == outSelIdx ? io_out_6_resp_bits_rdata : _GEN_65; // @[Decoupled.scala 40:37]
  wire  _GEN_77 = 3'h7 == outSelIdx ? io_out_7_req_ready : _GEN_66; // @[Decoupled.scala 40:37]
  wire  _GEN_78 = 3'h7 == outSelIdx ? io_out_7_req_valid : _GEN_67; // @[Decoupled.scala 40:37]
  wire [31:0] _GEN_79 = 3'h7 == outSelIdx ? io_out_7_req_bits_addr : _GEN_68; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_80 = 3'h7 == outSelIdx ? io_out_7_req_bits_size : _GEN_69; // @[Decoupled.scala 40:37]
  wire [3:0] _GEN_81 = 3'h7 == outSelIdx ? io_out_7_req_bits_cmd : _GEN_70; // @[Decoupled.scala 40:37]
  wire [7:0] _GEN_82 = 3'h7 == outSelIdx ? io_out_7_req_bits_wmask : _GEN_71; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_83 = 3'h7 == outSelIdx ? io_out_7_req_bits_wdata : _GEN_72; // @[Decoupled.scala 40:37]
  wire  _GEN_84 = 3'h7 == outSelIdx ? io_out_7_resp_ready : _GEN_73; // @[Decoupled.scala 40:37]
  wire  _GEN_85 = 3'h7 == outSelIdx ? io_out_7_resp_valid : _GEN_74; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_87 = 3'h7 == outSelIdx ? io_out_7_resp_bits_rdata : _GEN_76; // @[Decoupled.scala 40:37]
  wire  _T_30 = _GEN_77 & _GEN_78; // @[Decoupled.scala 40:37]
  wire  _T_31 = state == 2'h0; // @[Crossbar.scala 39:72]
  wire  _T_32 = _T_30 & _T_31; // @[Crossbar.scala 39:62]
  reg [2:0] outSelIdxResp; // @[Reg.scala 15:16]
  wire [7:0] _T_39 = {outSelVec_7,outSelVec_6,outSelVec_5,outSelVec_4,outSelVec_3,outSelVec_2,outSelVec_1,outSelVec_0}; // @[Crossbar.scala 41:54]
  wire  _T_40 = |_T_39; // @[Crossbar.scala 41:61]
  wire  _T_41 = ~_T_40; // @[Crossbar.scala 41:43]
  wire  reqInvalidAddr = io_in_req_valid & _T_41; // @[Crossbar.scala 41:40]
  wire  _T_59 = &_T_39; // @[Crossbar.scala 43:91]
  wire  _T_60 = io_in_req_valid & _T_59; // @[Crossbar.scala 43:71]
  wire  _T_61 = reqInvalidAddr | _T_60; // @[Crossbar.scala 43:51]
  reg [63:0] _T_64; // @[GTimer.scala 24:20]
  wire [63:0] _T_66 = _T_64 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_68 = ~reset; // @[Crossbar.scala 45:13]
  wire  _T_78 = ~_T_60; // @[Crossbar.scala 49:10]
  wire  _T_80 = _T_78 | reset; // @[Crossbar.scala 49:9]
  wire  _T_81 = ~_T_80; // @[Crossbar.scala 49:9]
  wire  _T_83 = io_in_req_valid & _T_31; // @[Crossbar.scala 54:42]
  wire  _T_106 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_108 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _GEN_109 = 3'h1 == outSelIdxResp ? io_out_1_resp_ready : io_out_0_resp_ready; // @[Decoupled.scala 40:37]
  wire  _GEN_110 = 3'h1 == outSelIdxResp ? io_out_1_resp_valid : io_out_0_resp_valid; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_112 = 3'h1 == outSelIdxResp ? io_out_1_resp_bits_rdata : io_out_0_resp_bits_rdata; // @[Decoupled.scala 40:37]
  wire  _GEN_120 = 3'h2 == outSelIdxResp ? io_out_2_resp_ready : _GEN_109; // @[Decoupled.scala 40:37]
  wire  _GEN_121 = 3'h2 == outSelIdxResp ? io_out_2_resp_valid : _GEN_110; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_123 = 3'h2 == outSelIdxResp ? io_out_2_resp_bits_rdata : _GEN_112; // @[Decoupled.scala 40:37]
  wire  _GEN_131 = 3'h3 == outSelIdxResp ? io_out_3_resp_ready : _GEN_120; // @[Decoupled.scala 40:37]
  wire  _GEN_132 = 3'h3 == outSelIdxResp ? io_out_3_resp_valid : _GEN_121; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_134 = 3'h3 == outSelIdxResp ? io_out_3_resp_bits_rdata : _GEN_123; // @[Decoupled.scala 40:37]
  wire  _GEN_142 = 3'h4 == outSelIdxResp ? io_out_4_resp_ready : _GEN_131; // @[Decoupled.scala 40:37]
  wire  _GEN_143 = 3'h4 == outSelIdxResp ? io_out_4_resp_valid : _GEN_132; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_145 = 3'h4 == outSelIdxResp ? io_out_4_resp_bits_rdata : _GEN_134; // @[Decoupled.scala 40:37]
  wire  _GEN_153 = 3'h5 == outSelIdxResp ? io_out_5_resp_ready : _GEN_142; // @[Decoupled.scala 40:37]
  wire  _GEN_154 = 3'h5 == outSelIdxResp ? io_out_5_resp_valid : _GEN_143; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_156 = 3'h5 == outSelIdxResp ? io_out_5_resp_bits_rdata : _GEN_145; // @[Decoupled.scala 40:37]
  wire  _GEN_164 = 3'h6 == outSelIdxResp ? io_out_6_resp_ready : _GEN_153; // @[Decoupled.scala 40:37]
  wire  _GEN_165 = 3'h6 == outSelIdxResp ? io_out_6_resp_valid : _GEN_154; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_167 = 3'h6 == outSelIdxResp ? io_out_6_resp_bits_rdata : _GEN_156; // @[Decoupled.scala 40:37]
  wire  _GEN_175 = 3'h7 == outSelIdxResp ? io_out_7_resp_ready : _GEN_164; // @[Decoupled.scala 40:37]
  wire  _GEN_176 = 3'h7 == outSelIdxResp ? io_out_7_resp_valid : _GEN_165; // @[Decoupled.scala 40:37]
  wire  _T_109 = _GEN_175 & _GEN_176; // @[Decoupled.scala 40:37]
  wire  _T_110 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_111 = io_in_resp_ready & io_in_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_113 = state == 2'h2; // @[Crossbar.scala 67:55]
  wire  _T_119 = _T_31 & io_in_req_valid; // @[Crossbar.scala 74:28]
  reg [63:0] _T_120; // @[GTimer.scala 24:20]
  wire [63:0] _T_122 = _T_120 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_126; // @[GTimer.scala 24:20]
  wire [63:0] _T_128 = _T_126 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_131 = _GEN_84 & _GEN_85; // @[Decoupled.scala 40:37]
  reg [63:0] _T_132; // @[GTimer.scala 24:20]
  wire [63:0] _T_134 = _T_132 + 64'h1; // @[GTimer.scala 25:12]
  reg [63:0] _T_138; // @[GTimer.scala 24:20]
  wire [63:0] _T_140 = _T_138 + 64'h1; // @[GTimer.scala 25:12]
  wire  _GEN_192 = _T_61 & DISPLAY_ENABLE; // @[Crossbar.scala 45:13]
  wire  _GEN_193 = DISPLAY_ENABLE & _T_119; // @[Crossbar.scala 75:13]
  wire  _GEN_194 = DISPLAY_ENABLE & _T_30; // @[Crossbar.scala 79:13]
  wire  _GEN_195 = DISPLAY_ENABLE & _T_131; // @[Crossbar.scala 82:13]
  wire  _GEN_196 = DISPLAY_ENABLE & _T_111; // @[Crossbar.scala 86:13]
  assign io_in_req_ready = _GEN_77 | reqInvalidAddr; // @[Crossbar.scala 71:19]
  assign io_in_resp_valid = _T_109 | _T_113; // @[Crossbar.scala 67:20]
  assign io_in_resp_bits_cmd = 4'h6; // @[Crossbar.scala 68:19]
  assign io_in_resp_bits_rdata = 3'h7 == outSelIdxResp ? io_out_7_resp_bits_rdata : _GEN_167; // @[Crossbar.scala 68:19]
  assign io_out_0_req_valid = outSelVec_0 & _T_83; // @[Crossbar.scala 54:17]
  assign io_out_0_req_bits_addr = io_in_req_bits_addr; // @[Crossbar.scala 53:16]
  assign io_out_0_req_bits_size = io_in_req_bits_size; // @[Crossbar.scala 53:16]
  assign io_out_0_req_bits_cmd = io_in_req_bits_cmd; // @[Crossbar.scala 53:16]
  assign io_out_0_req_bits_wmask = io_in_req_bits_wmask; // @[Crossbar.scala 53:16]
  assign io_out_0_req_bits_wdata = io_in_req_bits_wdata; // @[Crossbar.scala 53:16]
  assign io_out_0_resp_ready = 3'h0 == outSelIdxResp ? io_in_resp_ready : outSelVec_0; // @[Crossbar.scala 55:18 Crossbar.scala 70:25]
  assign io_out_1_req_valid = outSelVec_1 & _T_83; // @[Crossbar.scala 54:17]
  assign io_out_1_req_bits_addr = io_in_req_bits_addr; // @[Crossbar.scala 53:16]
  assign io_out_1_req_bits_size = io_in_req_bits_size; // @[Crossbar.scala 53:16]
  assign io_out_1_req_bits_cmd = io_in_req_bits_cmd; // @[Crossbar.scala 53:16]
  assign io_out_1_req_bits_wmask = io_in_req_bits_wmask; // @[Crossbar.scala 53:16]
  assign io_out_1_req_bits_wdata = io_in_req_bits_wdata; // @[Crossbar.scala 53:16]
  assign io_out_1_resp_ready = 3'h1 == outSelIdxResp ? io_in_resp_ready : outSelVec_1; // @[Crossbar.scala 55:18 Crossbar.scala 70:25]
  assign io_out_2_req_valid = outSelVec_2 & _T_83; // @[Crossbar.scala 54:17]
  assign io_out_2_req_bits_addr = io_in_req_bits_addr; // @[Crossbar.scala 53:16]
  assign io_out_2_req_bits_size = io_in_req_bits_size; // @[Crossbar.scala 53:16]
  assign io_out_2_req_bits_cmd = io_in_req_bits_cmd; // @[Crossbar.scala 53:16]
  assign io_out_2_req_bits_wmask = io_in_req_bits_wmask; // @[Crossbar.scala 53:16]
  assign io_out_2_req_bits_wdata = io_in_req_bits_wdata; // @[Crossbar.scala 53:16]
  assign io_out_2_resp_ready = 3'h2 == outSelIdxResp ? io_in_resp_ready : outSelVec_2; // @[Crossbar.scala 55:18 Crossbar.scala 70:25]
  assign io_out_3_req_valid = outSelVec_3 & _T_83; // @[Crossbar.scala 54:17]
  assign io_out_3_req_bits_addr = io_in_req_bits_addr; // @[Crossbar.scala 53:16]
  assign io_out_3_req_bits_size = io_in_req_bits_size; // @[Crossbar.scala 53:16]
  assign io_out_3_req_bits_cmd = io_in_req_bits_cmd; // @[Crossbar.scala 53:16]
  assign io_out_3_req_bits_wmask = io_in_req_bits_wmask; // @[Crossbar.scala 53:16]
  assign io_out_3_req_bits_wdata = io_in_req_bits_wdata; // @[Crossbar.scala 53:16]
  assign io_out_3_resp_ready = 3'h3 == outSelIdxResp ? io_in_resp_ready : outSelVec_3; // @[Crossbar.scala 55:18 Crossbar.scala 70:25]
  assign io_out_4_req_valid = outSelVec_4 & _T_83; // @[Crossbar.scala 54:17]
  assign io_out_4_req_bits_addr = io_in_req_bits_addr; // @[Crossbar.scala 53:16]
  assign io_out_4_req_bits_size = io_in_req_bits_size; // @[Crossbar.scala 53:16]
  assign io_out_4_req_bits_cmd = io_in_req_bits_cmd; // @[Crossbar.scala 53:16]
  assign io_out_4_req_bits_wmask = io_in_req_bits_wmask; // @[Crossbar.scala 53:16]
  assign io_out_4_req_bits_wdata = io_in_req_bits_wdata; // @[Crossbar.scala 53:16]
  assign io_out_4_resp_ready = 3'h4 == outSelIdxResp ? io_in_resp_ready : outSelVec_4; // @[Crossbar.scala 55:18 Crossbar.scala 70:25]
  assign io_out_5_req_valid = outSelVec_5 & _T_83; // @[Crossbar.scala 54:17]
  assign io_out_5_req_bits_addr = io_in_req_bits_addr; // @[Crossbar.scala 53:16]
  assign io_out_5_req_bits_size = io_in_req_bits_size; // @[Crossbar.scala 53:16]
  assign io_out_5_req_bits_cmd = io_in_req_bits_cmd; // @[Crossbar.scala 53:16]
  assign io_out_5_req_bits_wmask = io_in_req_bits_wmask; // @[Crossbar.scala 53:16]
  assign io_out_5_req_bits_wdata = io_in_req_bits_wdata; // @[Crossbar.scala 53:16]
  assign io_out_5_resp_ready = 3'h5 == outSelIdxResp ? io_in_resp_ready : outSelVec_5; // @[Crossbar.scala 55:18 Crossbar.scala 70:25]
  assign io_out_6_req_valid = outSelVec_6 & _T_83; // @[Crossbar.scala 54:17]
  assign io_out_6_req_bits_addr = io_in_req_bits_addr; // @[Crossbar.scala 53:16]
  assign io_out_6_req_bits_size = io_in_req_bits_size; // @[Crossbar.scala 53:16]
  assign io_out_6_req_bits_cmd = io_in_req_bits_cmd; // @[Crossbar.scala 53:16]
  assign io_out_6_req_bits_wmask = io_in_req_bits_wmask; // @[Crossbar.scala 53:16]
  assign io_out_6_req_bits_wdata = io_in_req_bits_wdata; // @[Crossbar.scala 53:16]
  assign io_out_6_resp_ready = 3'h6 == outSelIdxResp ? io_in_resp_ready : outSelVec_6; // @[Crossbar.scala 55:18 Crossbar.scala 70:25]
  assign io_out_7_req_valid = outSelVec_7 & _T_83; // @[Crossbar.scala 54:17]
  assign io_out_7_req_bits_addr = io_in_req_bits_addr; // @[Crossbar.scala 53:16]
  assign io_out_7_req_bits_size = io_in_req_bits_size; // @[Crossbar.scala 53:16]
  assign io_out_7_req_bits_cmd = io_in_req_bits_cmd; // @[Crossbar.scala 53:16]
  assign io_out_7_req_bits_wmask = io_in_req_bits_wmask; // @[Crossbar.scala 53:16]
  assign io_out_7_req_bits_wdata = io_in_req_bits_wdata; // @[Crossbar.scala 53:16]
  assign io_out_7_resp_ready = 3'h7 == outSelIdxResp ? io_in_resp_ready : outSelVec_7; // @[Crossbar.scala 55:18 Crossbar.scala 70:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  outSelIdxResp = _RAND_1[2:0];
  _RAND_2 = {2{`RANDOM}};
  _T_64 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  _T_120 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  _T_126 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  _T_132 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  _T_138 = _RAND_6[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else if (_T_106) begin
      if (reqInvalidAddr) begin
        state <= 2'h2;
      end else if (_T_30) begin
        state <= 2'h1;
      end
    end else if (_T_108) begin
      if (_T_109) begin
        state <= 2'h0;
      end
    end else if (_T_110) begin
      if (_T_111) begin
        state <= 2'h0;
      end
    end
    if (_T_32) begin
      if (outSelVec_0) begin
        outSelIdxResp <= 3'h0;
      end else if (outSelVec_1) begin
        outSelIdxResp <= 3'h1;
      end else if (outSelVec_2) begin
        outSelIdxResp <= 3'h2;
      end else if (outSelVec_3) begin
        outSelIdxResp <= 3'h3;
      end else if (outSelVec_4) begin
        outSelIdxResp <= 3'h4;
      end else if (outSelVec_5) begin
        outSelIdxResp <= 3'h5;
      end else if (outSelVec_6) begin
        outSelIdxResp <= 3'h6;
      end else begin
        outSelIdxResp <= 3'h7;
      end
    end
    if (reset) begin
      _T_64 <= 64'h0;
    end else begin
      _T_64 <= _T_66;
    end
    if (reset) begin
      _T_120 <= 64'h0;
    end else begin
      _T_120 <= _T_122;
    end
    if (reset) begin
      _T_126 <= 64'h0;
    end else begin
      _T_126 <= _T_128;
    end
    if (reset) begin
      _T_132 <= 64'h0;
    end else begin
      _T_132 <= _T_134;
    end
    if (reset) begin
      _T_138 <= 64'h0;
    end else begin
      _T_138 <= _T_140;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_192 & _T_68) begin
          $fwrite(32'h80000002,"crossbar access bad addr %x, time %d\n",io_in_req_bits_addr,_T_64); // @[Crossbar.scala 45:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_81) begin
          $fwrite(32'h80000002,"Assertion failed: address decode error, bad addr = 0x%x\n\n    at Crossbar.scala:49 assert(!(io.in.req.valid && outSelVec.asUInt.andR), \"address decode error, bad addr = 0x%%x\\n\", addr)\n",io_in_req_bits_addr); // @[Crossbar.scala 49:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_81) begin
          $fatal; // @[Crossbar.scala 49:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & _T_68) begin
          $fwrite(32'h80000002,"%d: xbar: in.req: addr = 0x%x, cmd = %d, size = %d, wmask = 0x%x, wdata = 0x%x\n",_T_120,io_in_req_bits_addr,io_in_req_bits_cmd,io_in_req_bits_size,io_in_req_bits_wmask,io_in_req_bits_wdata); // @[Crossbar.scala 75:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_194 & _T_68) begin
          $fwrite(32'h80000002,"%d: xbar: outSelIdx = %d, outSel.req: addr = 0x%x, cmd = %d, size = %d, wmask = 0x%x, wdata = 0x%x\n",_T_126,outSelIdx,_GEN_79,_GEN_81,_GEN_80,_GEN_82,_GEN_83); // @[Crossbar.scala 79:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_68) begin
          $fwrite(32'h80000002,"%d: xbar: outSelIdx= %d, outSel.resp: rdata = %x, cmd = %d\n",_T_132,outSelIdx,_GEN_87,4'h6); // @[Crossbar.scala 82:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_196 & _T_68) begin
          $fwrite(32'h80000002,"%d: xbar: in.resp: rdata = %x, cmd = %d\n",_T_138,io_in_resp_bits_rdata,io_in_resp_bits_cmd); // @[Crossbar.scala 86:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module AXI4UART(
  input         clock,
  input         reset,
  output        io_in_aw_ready,
  input         io_in_aw_valid,
  input  [31:0] io_in_aw_bits_addr,
  output        io_in_w_ready,
  input         io_in_w_valid,
  input  [63:0] io_in_w_bits_data,
  input  [7:0]  io_in_w_bits_strb,
  input         io_in_b_ready,
  output        io_in_b_valid,
  output        io_in_ar_ready,
  input         io_in_ar_valid,
  input  [31:0] io_in_ar_bits_addr,
  input         io_in_r_ready,
  output        io_in_r_valid,
  output [63:0] io_in_r_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  getcHelper_clk; // @[AXI4UART.scala 56:26]
  wire  getcHelper_getc; // @[AXI4UART.scala 56:26]
  wire [7:0] getcHelper_ch; // @[AXI4UART.scala 56:26]
  wire  _T_30 = io_in_ar_ready & io_in_ar_valid; // @[Decoupled.scala 40:37]
  wire  _T_31 = io_in_r_ready & io_in_r_valid; // @[Decoupled.scala 40:37]
  reg  r_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_31 ? 1'h0 : r_busy; // @[StopWatch.scala 26:19]
  wire  _GEN_1 = _T_30 | _GEN_0; // @[StopWatch.scala 27:20]
  wire  _T_33 = ~r_busy; // @[AXI4Slave.scala 71:32]
  reg  ren; // @[AXI4Slave.scala 73:17]
  wire  _T_42 = _T_30 | r_busy; // @[AXI4Slave.scala 74:52]
  wire  _T_43 = ren & _T_42; // @[AXI4Slave.scala 74:35]
  reg  _T_45; // @[StopWatch.scala 24:20]
  wire  _GEN_2 = _T_31 ? 1'h0 : _T_45; // @[StopWatch.scala 26:19]
  wire  _GEN_3 = _T_43 | _GEN_2; // @[StopWatch.scala 27:20]
  wire  _T_46 = io_in_aw_ready & io_in_aw_valid; // @[Decoupled.scala 40:37]
  wire  _T_47 = io_in_b_ready & io_in_b_valid; // @[Decoupled.scala 40:37]
  reg  w_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_4 = _T_47 ? 1'h0 : w_busy; // @[StopWatch.scala 26:19]
  wire  _GEN_5 = _T_46 | _GEN_4; // @[StopWatch.scala 27:20]
  wire  _T_50 = io_in_w_ready & io_in_w_valid; // @[Decoupled.scala 40:37]
  reg  _T_53; // @[StopWatch.scala 24:20]
  wire  _GEN_6 = _T_47 ? 1'h0 : _T_53; // @[StopWatch.scala 26:19]
  wire  _GEN_7 = _T_50 | _GEN_6; // @[StopWatch.scala 27:20]
  reg [31:0] txfifo; // @[AXI4UART.scala 52:19]
  reg [31:0] stat; // @[AXI4UART.scala 53:21]
  reg [31:0] ctrl; // @[AXI4UART.scala 54:21]
  wire  _T_55 = io_in_ar_bits_addr[3:0] == 4'h0; // @[AXI4UART.scala 58:37]
  wire [7:0] _T_61 = io_in_w_bits_strb >> io_in_aw_bits_addr[2:0]; // @[AXI4UART.scala 71:72]
  wire [7:0] _T_71 = _T_61[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_73 = _T_61[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_75 = _T_61[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_77 = _T_61[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_79 = _T_61[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_81 = _T_61[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_83 = _T_61[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_85 = _T_61[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_92 = {_T_85,_T_83,_T_81,_T_79,_T_77,_T_75,_T_73,_T_71}; // @[Cat.scala 29:58]
  wire  _T_93 = 4'h0 == io_in_ar_bits_addr[3:0]; // @[LookupTree.scala 24:34]
  wire  _T_94 = 4'h4 == io_in_ar_bits_addr[3:0]; // @[LookupTree.scala 24:34]
  wire  _T_95 = 4'h8 == io_in_ar_bits_addr[3:0]; // @[LookupTree.scala 24:34]
  wire  _T_96 = 4'hc == io_in_ar_bits_addr[3:0]; // @[LookupTree.scala 24:34]
  wire [7:0] _T_97 = _T_93 ? getcHelper_ch : 8'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_98 = _T_94 ? txfifo : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_99 = _T_95 ? stat : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_100 = _T_96 ? ctrl : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _GEN_11 = {{24'd0}, _T_97}; // @[Mux.scala 27:72]
  wire [31:0] _T_101 = _GEN_11 | _T_98; // @[Mux.scala 27:72]
  wire [31:0] _T_102 = _T_101 | _T_99; // @[Mux.scala 27:72]
  wire [31:0] _T_103 = _T_102 | _T_100; // @[Mux.scala 27:72]
  wire  _T_105 = io_in_aw_bits_addr[3:0] == 4'h4; // @[RegMap.scala 32:41]
  wire  _T_106 = _T_50 & _T_105; // @[RegMap.scala 32:32]
  wire [63:0] _T_107 = io_in_w_bits_data & _T_92; // @[BitUtils.scala 32:13]
  wire [63:0] _T_108 = ~_T_92; // @[BitUtils.scala 32:38]
  wire [63:0] _GEN_12 = {{32'd0}, txfifo}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_109 = _GEN_12 & _T_108; // @[BitUtils.scala 32:36]
  wire [63:0] _T_110 = _T_107 | _T_109; // @[BitUtils.scala 32:25]
  wire  _T_113 = ~reset; // @[AXI4UART.scala 60:37]
  wire [63:0] _GEN_8 = _T_106 ? _T_110 : {{32'd0}, txfifo}; // @[RegMap.scala 32:48]
  wire  _T_114 = io_in_aw_bits_addr[3:0] == 4'h8; // @[RegMap.scala 32:41]
  wire  _T_115 = _T_50 & _T_114; // @[RegMap.scala 32:32]
  wire [63:0] _GEN_13 = {{32'd0}, stat}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_118 = _GEN_13 & _T_108; // @[BitUtils.scala 32:36]
  wire [63:0] _T_119 = _T_107 | _T_118; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_9 = _T_115 ? _T_119 : {{32'd0}, stat}; // @[RegMap.scala 32:48]
  wire  _T_120 = io_in_aw_bits_addr[3:0] == 4'hc; // @[RegMap.scala 32:41]
  wire  _T_121 = _T_50 & _T_120; // @[RegMap.scala 32:32]
  wire [63:0] _GEN_14 = {{32'd0}, ctrl}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_124 = _GEN_14 & _T_108; // @[BitUtils.scala 32:36]
  wire [63:0] _T_125 = _T_107 | _T_124; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_10 = _T_121 ? _T_125 : {{32'd0}, ctrl}; // @[RegMap.scala 32:48]
  UARTGetc getcHelper ( // @[AXI4UART.scala 56:26]
    .clk(getcHelper_clk),
    .getc(getcHelper_getc),
    .ch(getcHelper_ch)
  );
  assign io_in_aw_ready = ~w_busy; // @[AXI4Slave.scala 94:15]
  assign io_in_w_ready = io_in_aw_valid | w_busy; // @[AXI4Slave.scala 95:15]
  assign io_in_b_valid = _T_53; // @[AXI4Slave.scala 97:14]
  assign io_in_ar_ready = io_in_r_ready | _T_33; // @[AXI4Slave.scala 71:15]
  assign io_in_r_valid = _T_45; // @[AXI4Slave.scala 74:14]
  assign io_in_r_bits_data = {{32'd0}, _T_103}; // @[RegMap.scala 30:11]
  assign getcHelper_clk = clock; // @[AXI4UART.scala 57:21]
  assign getcHelper_getc = _T_55 & ren; // @[AXI4UART.scala 58:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ren = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _T_45 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_53 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  txfifo = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  stat = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  ctrl = _RAND_7[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      r_busy <= 1'h0;
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin
      ren <= 1'h0;
    end else begin
      ren <= _T_30;
    end
    if (reset) begin
      _T_45 <= 1'h0;
    end else begin
      _T_45 <= _GEN_3;
    end
    if (reset) begin
      w_busy <= 1'h0;
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin
      _T_53 <= 1'h0;
    end else begin
      _T_53 <= _GEN_7;
    end
    txfifo <= _GEN_8[31:0];
    if (reset) begin
      stat <= 32'h1;
    end else begin
      stat <= _GEN_9[31:0];
    end
    if (reset) begin
      ctrl <= 32'h0;
    end else begin
      ctrl <= _GEN_10[31:0];
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_106 & _T_113) begin
          $fwrite(32'h80000002,"%c",_T_110[7:0]); // @[AXI4UART.scala 60:37]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module VGACtrl(
  input         clock,
  input         reset,
  output        io_in_aw_ready,
  input         io_in_aw_valid,
  output        io_in_w_ready,
  input         io_in_w_valid,
  input         io_in_b_ready,
  output        io_in_b_valid,
  output        io_in_ar_ready,
  input         io_in_ar_valid,
  input  [31:0] io_in_ar_bits_addr,
  input         io_in_r_ready,
  output        io_in_r_valid,
  output [63:0] io_in_r_bits_data,
  output        io_extra_sync
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  _T_30 = io_in_ar_ready & io_in_ar_valid; // @[Decoupled.scala 40:37]
  wire  _T_31 = io_in_r_ready & io_in_r_valid; // @[Decoupled.scala 40:37]
  reg  r_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_31 ? 1'h0 : r_busy; // @[StopWatch.scala 26:19]
  wire  _GEN_1 = _T_30 | _GEN_0; // @[StopWatch.scala 27:20]
  wire  _T_33 = ~r_busy; // @[AXI4Slave.scala 71:32]
  reg  ren; // @[AXI4Slave.scala 73:17]
  wire  _T_42 = _T_30 | r_busy; // @[AXI4Slave.scala 74:52]
  wire  _T_43 = ren & _T_42; // @[AXI4Slave.scala 74:35]
  reg  _T_45; // @[StopWatch.scala 24:20]
  wire  _GEN_2 = _T_31 ? 1'h0 : _T_45; // @[StopWatch.scala 26:19]
  wire  _GEN_3 = _T_43 | _GEN_2; // @[StopWatch.scala 27:20]
  wire  _T_46 = io_in_aw_ready & io_in_aw_valid; // @[Decoupled.scala 40:37]
  wire  _T_47 = io_in_b_ready & io_in_b_valid; // @[Decoupled.scala 40:37]
  reg  w_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_4 = _T_47 ? 1'h0 : w_busy; // @[StopWatch.scala 26:19]
  wire  _GEN_5 = _T_46 | _GEN_4; // @[StopWatch.scala 27:20]
  wire  _T_50 = io_in_w_ready & io_in_w_valid; // @[Decoupled.scala 40:37]
  reg  _T_53; // @[StopWatch.scala 24:20]
  wire  _GEN_6 = _T_47 ? 1'h0 : _T_53; // @[StopWatch.scala 26:19]
  wire  _GEN_7 = _T_50 | _GEN_6; // @[StopWatch.scala 27:20]
  wire  _T_88 = 4'h0 == io_in_ar_bits_addr[3:0]; // @[LookupTree.scala 24:34]
  wire  _T_89 = 4'h4 == io_in_ar_bits_addr[3:0]; // @[LookupTree.scala 24:34]
  wire [31:0] _T_90 = _T_88 ? 32'h190012c : 32'h0; // @[Mux.scala 27:72]
  wire  _T_91 = _T_89 & _T_46; // @[Mux.scala 27:72]
  wire [31:0] _GEN_8 = {{31'd0}, _T_91}; // @[Mux.scala 27:72]
  wire [31:0] _T_92 = _T_90 | _GEN_8; // @[Mux.scala 27:72]
  assign io_in_aw_ready = ~w_busy; // @[AXI4Slave.scala 94:15]
  assign io_in_w_ready = io_in_aw_valid | w_busy; // @[AXI4Slave.scala 95:15]
  assign io_in_b_valid = _T_53; // @[AXI4Slave.scala 97:14]
  assign io_in_ar_ready = io_in_r_ready | _T_33; // @[AXI4Slave.scala 71:15]
  assign io_in_r_valid = _T_45; // @[AXI4Slave.scala 74:14]
  assign io_in_r_bits_data = {{32'd0}, _T_92}; // @[RegMap.scala 30:11]
  assign io_extra_sync = io_in_aw_ready & io_in_aw_valid; // @[AXI4VGA.scala 83:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ren = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _T_45 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_53 = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      r_busy <= 1'h0;
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin
      ren <= 1'h0;
    end else begin
      ren <= _T_30;
    end
    if (reset) begin
      _T_45 <= 1'h0;
    end else begin
      _T_45 <= _GEN_3;
    end
    if (reset) begin
      w_busy <= 1'h0;
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin
      _T_53 <= 1'h0;
    end else begin
      _T_53 <= _GEN_7;
    end
  end
endmodule
module AXI4RAM_1(
  input         clock,
  input         reset,
  output        io_in_aw_ready,
  input         io_in_aw_valid,
  input  [31:0] io_in_aw_bits_addr,
  output        io_in_w_ready,
  input         io_in_w_valid,
  input  [63:0] io_in_w_bits_data,
  input  [7:0]  io_in_w_bits_strb,
  input         io_in_b_ready,
  output        io_in_b_valid,
  output        io_in_ar_ready,
  input         io_in_ar_valid,
  input  [31:0] io_in_ar_bits_addr,
  input         io_in_r_ready,
  output        io_in_r_valid,
  output [63:0] io_in_r_bits_data
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [63:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] _T_62_0 [0:59999]; // @[AXI4RAM.scala 61:18]
  wire [7:0] _T_62_0__T_85_data; // @[AXI4RAM.scala 61:18]
  wire [15:0] _T_62_0__T_85_addr; // @[AXI4RAM.scala 61:18]
  wire [7:0] _T_62_0__T_82_data; // @[AXI4RAM.scala 61:18]
  wire [15:0] _T_62_0__T_82_addr; // @[AXI4RAM.scala 61:18]
  wire  _T_62_0__T_82_mask; // @[AXI4RAM.scala 61:18]
  wire  _T_62_0__T_82_en; // @[AXI4RAM.scala 61:18]
  reg [7:0] _T_62_1 [0:59999]; // @[AXI4RAM.scala 61:18]
  wire [7:0] _T_62_1__T_85_data; // @[AXI4RAM.scala 61:18]
  wire [15:0] _T_62_1__T_85_addr; // @[AXI4RAM.scala 61:18]
  wire [7:0] _T_62_1__T_82_data; // @[AXI4RAM.scala 61:18]
  wire [15:0] _T_62_1__T_82_addr; // @[AXI4RAM.scala 61:18]
  wire  _T_62_1__T_82_mask; // @[AXI4RAM.scala 61:18]
  wire  _T_62_1__T_82_en; // @[AXI4RAM.scala 61:18]
  reg [7:0] _T_62_2 [0:59999]; // @[AXI4RAM.scala 61:18]
  wire [7:0] _T_62_2__T_85_data; // @[AXI4RAM.scala 61:18]
  wire [15:0] _T_62_2__T_85_addr; // @[AXI4RAM.scala 61:18]
  wire [7:0] _T_62_2__T_82_data; // @[AXI4RAM.scala 61:18]
  wire [15:0] _T_62_2__T_82_addr; // @[AXI4RAM.scala 61:18]
  wire  _T_62_2__T_82_mask; // @[AXI4RAM.scala 61:18]
  wire  _T_62_2__T_82_en; // @[AXI4RAM.scala 61:18]
  reg [7:0] _T_62_3 [0:59999]; // @[AXI4RAM.scala 61:18]
  wire [7:0] _T_62_3__T_85_data; // @[AXI4RAM.scala 61:18]
  wire [15:0] _T_62_3__T_85_addr; // @[AXI4RAM.scala 61:18]
  wire [7:0] _T_62_3__T_82_data; // @[AXI4RAM.scala 61:18]
  wire [15:0] _T_62_3__T_82_addr; // @[AXI4RAM.scala 61:18]
  wire  _T_62_3__T_82_mask; // @[AXI4RAM.scala 61:18]
  wire  _T_62_3__T_82_en; // @[AXI4RAM.scala 61:18]
  reg [7:0] _T_62_4 [0:59999]; // @[AXI4RAM.scala 61:18]
  wire [7:0] _T_62_4__T_85_data; // @[AXI4RAM.scala 61:18]
  wire [15:0] _T_62_4__T_85_addr; // @[AXI4RAM.scala 61:18]
  wire [7:0] _T_62_4__T_82_data; // @[AXI4RAM.scala 61:18]
  wire [15:0] _T_62_4__T_82_addr; // @[AXI4RAM.scala 61:18]
  wire  _T_62_4__T_82_mask; // @[AXI4RAM.scala 61:18]
  wire  _T_62_4__T_82_en; // @[AXI4RAM.scala 61:18]
  reg [7:0] _T_62_5 [0:59999]; // @[AXI4RAM.scala 61:18]
  wire [7:0] _T_62_5__T_85_data; // @[AXI4RAM.scala 61:18]
  wire [15:0] _T_62_5__T_85_addr; // @[AXI4RAM.scala 61:18]
  wire [7:0] _T_62_5__T_82_data; // @[AXI4RAM.scala 61:18]
  wire [15:0] _T_62_5__T_82_addr; // @[AXI4RAM.scala 61:18]
  wire  _T_62_5__T_82_mask; // @[AXI4RAM.scala 61:18]
  wire  _T_62_5__T_82_en; // @[AXI4RAM.scala 61:18]
  reg [7:0] _T_62_6 [0:59999]; // @[AXI4RAM.scala 61:18]
  wire [7:0] _T_62_6__T_85_data; // @[AXI4RAM.scala 61:18]
  wire [15:0] _T_62_6__T_85_addr; // @[AXI4RAM.scala 61:18]
  wire [7:0] _T_62_6__T_82_data; // @[AXI4RAM.scala 61:18]
  wire [15:0] _T_62_6__T_82_addr; // @[AXI4RAM.scala 61:18]
  wire  _T_62_6__T_82_mask; // @[AXI4RAM.scala 61:18]
  wire  _T_62_6__T_82_en; // @[AXI4RAM.scala 61:18]
  reg [7:0] _T_62_7 [0:59999]; // @[AXI4RAM.scala 61:18]
  wire [7:0] _T_62_7__T_85_data; // @[AXI4RAM.scala 61:18]
  wire [15:0] _T_62_7__T_85_addr; // @[AXI4RAM.scala 61:18]
  wire [7:0] _T_62_7__T_82_data; // @[AXI4RAM.scala 61:18]
  wire [15:0] _T_62_7__T_82_addr; // @[AXI4RAM.scala 61:18]
  wire  _T_62_7__T_82_mask; // @[AXI4RAM.scala 61:18]
  wire  _T_62_7__T_82_en; // @[AXI4RAM.scala 61:18]
  wire  _T_30 = io_in_ar_ready & io_in_ar_valid; // @[Decoupled.scala 40:37]
  reg  r_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = io_in_r_valid ? 1'h0 : r_busy; // @[StopWatch.scala 26:19]
  wire  _GEN_1 = _T_30 | _GEN_0; // @[StopWatch.scala 27:20]
  reg  ren; // @[AXI4Slave.scala 73:17]
  wire  _T_42 = _T_30 | r_busy; // @[AXI4Slave.scala 74:52]
  wire  _T_43 = ren & _T_42; // @[AXI4Slave.scala 74:35]
  reg  _T_45; // @[StopWatch.scala 24:20]
  wire  _GEN_2 = io_in_r_valid ? 1'h0 : _T_45; // @[StopWatch.scala 26:19]
  wire  _GEN_3 = _T_43 | _GEN_2; // @[StopWatch.scala 27:20]
  wire  _T_46 = io_in_aw_ready & io_in_aw_valid; // @[Decoupled.scala 40:37]
  wire  _T_47 = io_in_b_ready & io_in_b_valid; // @[Decoupled.scala 40:37]
  reg  w_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_4 = _T_47 ? 1'h0 : w_busy; // @[StopWatch.scala 26:19]
  wire  _GEN_5 = _T_46 | _GEN_4; // @[StopWatch.scala 27:20]
  wire  _T_50 = io_in_w_ready & io_in_w_valid; // @[Decoupled.scala 40:37]
  reg  _T_53; // @[StopWatch.scala 24:20]
  wire  _GEN_6 = _T_47 ? 1'h0 : _T_53; // @[StopWatch.scala 26:19]
  wire  _GEN_7 = _T_50 | _GEN_6; // @[StopWatch.scala 27:20]
  wire [31:0] _T_54 = io_in_aw_bits_addr & 32'h7ffff; // @[AXI4RAM.scala 44:33]
  wire [29:0] _T_56 = {{1'd0}, _T_54[31:3]}; // @[AXI4RAM.scala 47:27]
  wire [28:0] wIdx = _T_56[28:0]; // @[AXI4RAM.scala 47:27]
  wire [31:0] _T_57 = io_in_ar_bits_addr & 32'h7ffff; // @[AXI4RAM.scala 44:33]
  wire [29:0] _T_59 = {{1'd0}, _T_57[31:3]}; // @[AXI4RAM.scala 48:27]
  wire [28:0] rIdx = _T_59[28:0]; // @[AXI4RAM.scala 48:27]
  wire  _T_61 = wIdx < 29'hea60; // @[AXI4RAM.scala 45:32]
  wire [63:0] rdata = {_T_62_7__T_85_data,_T_62_6__T_85_data,_T_62_5__T_85_data,_T_62_4__T_85_data,_T_62_3__T_85_data,_T_62_2__T_85_data,_T_62_1__T_85_data,_T_62_0__T_85_data}; // @[Cat.scala 29:58]
  reg [63:0] _T_92; // @[Reg.scala 15:16]
  assign _T_62_0__T_85_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_62_0__T_85_data = _T_62_0[_T_62_0__T_85_addr]; // @[AXI4RAM.scala 61:18]
  `else
  assign _T_62_0__T_85_data = _T_62_0__T_85_addr >= 16'hea60 ? _RAND_1[7:0] : _T_62_0[_T_62_0__T_85_addr]; // @[AXI4RAM.scala 61:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_62_0__T_82_data = io_in_w_bits_data[7:0];
  assign _T_62_0__T_82_addr = wIdx[15:0];
  assign _T_62_0__T_82_mask = io_in_w_bits_strb[0];
  assign _T_62_0__T_82_en = _T_50 & _T_61;
  assign _T_62_1__T_85_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_62_1__T_85_data = _T_62_1[_T_62_1__T_85_addr]; // @[AXI4RAM.scala 61:18]
  `else
  assign _T_62_1__T_85_data = _T_62_1__T_85_addr >= 16'hea60 ? _RAND_3[7:0] : _T_62_1[_T_62_1__T_85_addr]; // @[AXI4RAM.scala 61:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_62_1__T_82_data = io_in_w_bits_data[15:8];
  assign _T_62_1__T_82_addr = wIdx[15:0];
  assign _T_62_1__T_82_mask = io_in_w_bits_strb[1];
  assign _T_62_1__T_82_en = _T_50 & _T_61;
  assign _T_62_2__T_85_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_62_2__T_85_data = _T_62_2[_T_62_2__T_85_addr]; // @[AXI4RAM.scala 61:18]
  `else
  assign _T_62_2__T_85_data = _T_62_2__T_85_addr >= 16'hea60 ? _RAND_5[7:0] : _T_62_2[_T_62_2__T_85_addr]; // @[AXI4RAM.scala 61:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_62_2__T_82_data = io_in_w_bits_data[23:16];
  assign _T_62_2__T_82_addr = wIdx[15:0];
  assign _T_62_2__T_82_mask = io_in_w_bits_strb[2];
  assign _T_62_2__T_82_en = _T_50 & _T_61;
  assign _T_62_3__T_85_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_62_3__T_85_data = _T_62_3[_T_62_3__T_85_addr]; // @[AXI4RAM.scala 61:18]
  `else
  assign _T_62_3__T_85_data = _T_62_3__T_85_addr >= 16'hea60 ? _RAND_7[7:0] : _T_62_3[_T_62_3__T_85_addr]; // @[AXI4RAM.scala 61:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_62_3__T_82_data = io_in_w_bits_data[31:24];
  assign _T_62_3__T_82_addr = wIdx[15:0];
  assign _T_62_3__T_82_mask = io_in_w_bits_strb[3];
  assign _T_62_3__T_82_en = _T_50 & _T_61;
  assign _T_62_4__T_85_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_62_4__T_85_data = _T_62_4[_T_62_4__T_85_addr]; // @[AXI4RAM.scala 61:18]
  `else
  assign _T_62_4__T_85_data = _T_62_4__T_85_addr >= 16'hea60 ? _RAND_9[7:0] : _T_62_4[_T_62_4__T_85_addr]; // @[AXI4RAM.scala 61:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_62_4__T_82_data = io_in_w_bits_data[39:32];
  assign _T_62_4__T_82_addr = wIdx[15:0];
  assign _T_62_4__T_82_mask = io_in_w_bits_strb[4];
  assign _T_62_4__T_82_en = _T_50 & _T_61;
  assign _T_62_5__T_85_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_62_5__T_85_data = _T_62_5[_T_62_5__T_85_addr]; // @[AXI4RAM.scala 61:18]
  `else
  assign _T_62_5__T_85_data = _T_62_5__T_85_addr >= 16'hea60 ? _RAND_11[7:0] : _T_62_5[_T_62_5__T_85_addr]; // @[AXI4RAM.scala 61:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_62_5__T_82_data = io_in_w_bits_data[47:40];
  assign _T_62_5__T_82_addr = wIdx[15:0];
  assign _T_62_5__T_82_mask = io_in_w_bits_strb[5];
  assign _T_62_5__T_82_en = _T_50 & _T_61;
  assign _T_62_6__T_85_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_62_6__T_85_data = _T_62_6[_T_62_6__T_85_addr]; // @[AXI4RAM.scala 61:18]
  `else
  assign _T_62_6__T_85_data = _T_62_6__T_85_addr >= 16'hea60 ? _RAND_13[7:0] : _T_62_6[_T_62_6__T_85_addr]; // @[AXI4RAM.scala 61:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_62_6__T_82_data = io_in_w_bits_data[55:48];
  assign _T_62_6__T_82_addr = wIdx[15:0];
  assign _T_62_6__T_82_mask = io_in_w_bits_strb[6];
  assign _T_62_6__T_82_en = _T_50 & _T_61;
  assign _T_62_7__T_85_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_62_7__T_85_data = _T_62_7[_T_62_7__T_85_addr]; // @[AXI4RAM.scala 61:18]
  `else
  assign _T_62_7__T_85_data = _T_62_7__T_85_addr >= 16'hea60 ? _RAND_15[7:0] : _T_62_7[_T_62_7__T_85_addr]; // @[AXI4RAM.scala 61:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_62_7__T_82_data = io_in_w_bits_data[63:56];
  assign _T_62_7__T_82_addr = wIdx[15:0];
  assign _T_62_7__T_82_mask = io_in_w_bits_strb[7];
  assign _T_62_7__T_82_en = _T_50 & _T_61;
  assign io_in_aw_ready = ~w_busy; // @[AXI4Slave.scala 94:15]
  assign io_in_w_ready = io_in_aw_valid | w_busy; // @[AXI4Slave.scala 95:15]
  assign io_in_b_valid = _T_53; // @[AXI4Slave.scala 97:14]
  assign io_in_ar_ready = 1'h1; // @[AXI4Slave.scala 71:15]
  assign io_in_r_valid = _T_45; // @[AXI4Slave.scala 74:14]
  assign io_in_r_bits_data = _T_92; // @[AXI4RAM.scala 69:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_3 = {1{`RANDOM}};
  _RAND_5 = {1{`RANDOM}};
  _RAND_7 = {1{`RANDOM}};
  _RAND_9 = {1{`RANDOM}};
  _RAND_11 = {1{`RANDOM}};
  _RAND_13 = {1{`RANDOM}};
  _RAND_15 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    _T_62_0[initvar] = _RAND_0[7:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    _T_62_1[initvar] = _RAND_2[7:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    _T_62_2[initvar] = _RAND_4[7:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    _T_62_3[initvar] = _RAND_6[7:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    _T_62_4[initvar] = _RAND_8[7:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    _T_62_5[initvar] = _RAND_10[7:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    _T_62_6[initvar] = _RAND_12[7:0];
  _RAND_14 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    _T_62_7[initvar] = _RAND_14[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  r_busy = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  ren = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  _T_45 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  w_busy = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  _T_53 = _RAND_20[0:0];
  _RAND_21 = {2{`RANDOM}};
  _T_92 = _RAND_21[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_62_0__T_82_en & _T_62_0__T_82_mask) begin
      _T_62_0[_T_62_0__T_82_addr] <= _T_62_0__T_82_data; // @[AXI4RAM.scala 61:18]
    end
    if(_T_62_1__T_82_en & _T_62_1__T_82_mask) begin
      _T_62_1[_T_62_1__T_82_addr] <= _T_62_1__T_82_data; // @[AXI4RAM.scala 61:18]
    end
    if(_T_62_2__T_82_en & _T_62_2__T_82_mask) begin
      _T_62_2[_T_62_2__T_82_addr] <= _T_62_2__T_82_data; // @[AXI4RAM.scala 61:18]
    end
    if(_T_62_3__T_82_en & _T_62_3__T_82_mask) begin
      _T_62_3[_T_62_3__T_82_addr] <= _T_62_3__T_82_data; // @[AXI4RAM.scala 61:18]
    end
    if(_T_62_4__T_82_en & _T_62_4__T_82_mask) begin
      _T_62_4[_T_62_4__T_82_addr] <= _T_62_4__T_82_data; // @[AXI4RAM.scala 61:18]
    end
    if(_T_62_5__T_82_en & _T_62_5__T_82_mask) begin
      _T_62_5[_T_62_5__T_82_addr] <= _T_62_5__T_82_data; // @[AXI4RAM.scala 61:18]
    end
    if(_T_62_6__T_82_en & _T_62_6__T_82_mask) begin
      _T_62_6[_T_62_6__T_82_addr] <= _T_62_6__T_82_data; // @[AXI4RAM.scala 61:18]
    end
    if(_T_62_7__T_82_en & _T_62_7__T_82_mask) begin
      _T_62_7[_T_62_7__T_82_addr] <= _T_62_7__T_82_data; // @[AXI4RAM.scala 61:18]
    end
    if (reset) begin
      r_busy <= 1'h0;
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin
      ren <= 1'h0;
    end else begin
      ren <= _T_30;
    end
    if (reset) begin
      _T_45 <= 1'h0;
    end else begin
      _T_45 <= _GEN_3;
    end
    if (reset) begin
      w_busy <= 1'h0;
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin
      _T_53 <= 1'h0;
    end else begin
      _T_53 <= _GEN_7;
    end
    if (ren) begin
      _T_92 <= rdata;
    end
  end
endmodule
module AXI4VGA(
  input         clock,
  input         reset,
  output        io_in_fb_aw_ready,
  input         io_in_fb_aw_valid,
  input  [31:0] io_in_fb_aw_bits_addr,
  output        io_in_fb_w_ready,
  input         io_in_fb_w_valid,
  input  [63:0] io_in_fb_w_bits_data,
  input  [7:0]  io_in_fb_w_bits_strb,
  input         io_in_fb_b_ready,
  output        io_in_fb_b_valid,
  output        io_in_fb_ar_ready,
  input         io_in_fb_ar_valid,
  input         io_in_fb_r_ready,
  output        io_in_fb_r_valid,
  output        io_in_ctrl_aw_ready,
  input         io_in_ctrl_aw_valid,
  output        io_in_ctrl_w_ready,
  input         io_in_ctrl_w_valid,
  input         io_in_ctrl_b_ready,
  output        io_in_ctrl_b_valid,
  output        io_in_ctrl_ar_ready,
  input         io_in_ctrl_ar_valid,
  input  [31:0] io_in_ctrl_ar_bits_addr,
  input         io_in_ctrl_r_ready,
  output        io_in_ctrl_r_valid,
  output [63:0] io_in_ctrl_r_bits_data,
  output        io_vga_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  ctrl_clock; // @[AXI4VGA.scala 125:20]
  wire  ctrl_reset; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_aw_ready; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_aw_valid; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_w_ready; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_w_valid; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_b_ready; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_b_valid; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_ar_ready; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_ar_valid; // @[AXI4VGA.scala 125:20]
  wire [31:0] ctrl_io_in_ar_bits_addr; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_r_ready; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_r_valid; // @[AXI4VGA.scala 125:20]
  wire [63:0] ctrl_io_in_r_bits_data; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_extra_sync; // @[AXI4VGA.scala 125:20]
  wire  fb_clock; // @[AXI4VGA.scala 127:18]
  wire  fb_reset; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_aw_ready; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_aw_valid; // @[AXI4VGA.scala 127:18]
  wire [31:0] fb_io_in_aw_bits_addr; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_w_ready; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_w_valid; // @[AXI4VGA.scala 127:18]
  wire [63:0] fb_io_in_w_bits_data; // @[AXI4VGA.scala 127:18]
  wire [7:0] fb_io_in_w_bits_strb; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_b_ready; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_b_valid; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_ar_ready; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_ar_valid; // @[AXI4VGA.scala 127:18]
  wire [31:0] fb_io_in_ar_bits_addr; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_r_ready; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_r_valid; // @[AXI4VGA.scala 127:18]
  wire [63:0] fb_io_in_r_bits_data; // @[AXI4VGA.scala 127:18]
  wire  FBHelper_clk; // @[AXI4VGA.scala 171:26]
  wire  FBHelper_valid; // @[AXI4VGA.scala 171:26]
  wire [31:0] FBHelper_pixel; // @[AXI4VGA.scala 171:26]
  wire  FBHelper_sync; // @[AXI4VGA.scala 171:26]
  wire  _T = io_in_fb_ar_ready & io_in_fb_ar_valid; // @[Decoupled.scala 40:37]
  wire  _T_1 = io_in_fb_r_ready & io_in_fb_r_valid; // @[Decoupled.scala 40:37]
  reg  _T_2; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_1 ? 1'h0 : _T_2; // @[StopWatch.scala 26:19]
  wire  _GEN_1 = _T | _GEN_0; // @[StopWatch.scala 27:20]
  reg [10:0] hCounter; // @[Counter.scala 29:33]
  wire  hFinish = hCounter == 11'h41f; // @[Counter.scala 38:24]
  wire [10:0] _T_5 = hCounter + 11'h1; // @[Counter.scala 39:22]
  reg [9:0] vCounter; // @[Counter.scala 29:33]
  wire  _T_6 = vCounter == 10'h273; // @[Counter.scala 38:24]
  wire [9:0] _T_8 = vCounter + 10'h1; // @[Counter.scala 39:22]
  wire  _T_11 = hCounter >= 11'ha8; // @[AXI4VGA.scala 138:51]
  wire  _T_12 = hCounter < 11'h3c8; // @[AXI4VGA.scala 138:69]
  wire  hInRange = _T_11 & _T_12; // @[AXI4VGA.scala 138:63]
  wire  _T_13 = vCounter >= 10'h5; // @[AXI4VGA.scala 138:51]
  wire  _T_14 = vCounter < 10'h25d; // @[AXI4VGA.scala 138:69]
  wire  vInRange = _T_13 & _T_14; // @[AXI4VGA.scala 138:63]
  wire  hCounterIsOdd = hCounter[0]; // @[AXI4VGA.scala 150:31]
  wire  hCounterIs2 = hCounter[1:0] == 2'h2; // @[AXI4VGA.scala 151:35]
  wire  vCounterIsOdd = vCounter[0]; // @[AXI4VGA.scala 152:31]
  wire  _T_17 = hCounter >= 11'ha7; // @[AXI4VGA.scala 138:51]
  wire  _T_18 = hCounter < 11'h3c7; // @[AXI4VGA.scala 138:69]
  wire  _T_19 = _T_17 & _T_18; // @[AXI4VGA.scala 138:63]
  wire  _T_20 = _T_19 & vInRange; // @[AXI4VGA.scala 155:66]
  wire  nextPixel = _T_20 & hCounterIsOdd; // @[AXI4VGA.scala 155:78]
  wire  _T_21 = ~vCounterIsOdd; // @[AXI4VGA.scala 156:44]
  wire  _T_22 = nextPixel & _T_21; // @[AXI4VGA.scala 156:41]
  reg [16:0] fbPixelAddrV0; // @[Counter.scala 29:33]
  wire  _T_24 = fbPixelAddrV0 == 17'h1d4bf; // @[Counter.scala 38:24]
  wire [16:0] _T_26 = fbPixelAddrV0 + 17'h1; // @[Counter.scala 39:22]
  wire  _T_27 = nextPixel & vCounterIsOdd; // @[AXI4VGA.scala 157:41]
  reg [16:0] fbPixelAddrV1; // @[Counter.scala 29:33]
  wire  _T_29 = fbPixelAddrV1 == 17'h1d4bf; // @[Counter.scala 38:24]
  wire [16:0] _T_31 = fbPixelAddrV1 + 17'h1; // @[Counter.scala 39:22]
  wire [16:0] _T_32 = vCounterIsOdd ? fbPixelAddrV1 : fbPixelAddrV0; // @[AXI4VGA.scala 161:35]
  wire [18:0] _T_33 = {_T_32,2'h0}; // @[Cat.scala 29:58]
  reg  _T_34; // @[AXI4VGA.scala 162:31]
  wire  _T_36 = fb_io_in_r_ready & fb_io_in_r_valid; // @[Decoupled.scala 40:37]
  reg [63:0] _T_38; // @[Reg.scala 27:20]
  wire [63:0] _GEN_14 = _T_36 ? fb_io_in_r_bits_data : _T_38; // @[Reg.scala 28:19]
  VGACtrl ctrl ( // @[AXI4VGA.scala 125:20]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_in_aw_ready(ctrl_io_in_aw_ready),
    .io_in_aw_valid(ctrl_io_in_aw_valid),
    .io_in_w_ready(ctrl_io_in_w_ready),
    .io_in_w_valid(ctrl_io_in_w_valid),
    .io_in_b_ready(ctrl_io_in_b_ready),
    .io_in_b_valid(ctrl_io_in_b_valid),
    .io_in_ar_ready(ctrl_io_in_ar_ready),
    .io_in_ar_valid(ctrl_io_in_ar_valid),
    .io_in_ar_bits_addr(ctrl_io_in_ar_bits_addr),
    .io_in_r_ready(ctrl_io_in_r_ready),
    .io_in_r_valid(ctrl_io_in_r_valid),
    .io_in_r_bits_data(ctrl_io_in_r_bits_data),
    .io_extra_sync(ctrl_io_extra_sync)
  );
  AXI4RAM_1 fb ( // @[AXI4VGA.scala 127:18]
    .clock(fb_clock),
    .reset(fb_reset),
    .io_in_aw_ready(fb_io_in_aw_ready),
    .io_in_aw_valid(fb_io_in_aw_valid),
    .io_in_aw_bits_addr(fb_io_in_aw_bits_addr),
    .io_in_w_ready(fb_io_in_w_ready),
    .io_in_w_valid(fb_io_in_w_valid),
    .io_in_w_bits_data(fb_io_in_w_bits_data),
    .io_in_w_bits_strb(fb_io_in_w_bits_strb),
    .io_in_b_ready(fb_io_in_b_ready),
    .io_in_b_valid(fb_io_in_b_valid),
    .io_in_ar_ready(fb_io_in_ar_ready),
    .io_in_ar_valid(fb_io_in_ar_valid),
    .io_in_ar_bits_addr(fb_io_in_ar_bits_addr),
    .io_in_r_ready(fb_io_in_r_ready),
    .io_in_r_valid(fb_io_in_r_valid),
    .io_in_r_bits_data(fb_io_in_r_bits_data)
  );
  FBHelper FBHelper ( // @[AXI4VGA.scala 171:26]
    .clk(FBHelper_clk),
    .valid(FBHelper_valid),
    .pixel(FBHelper_pixel),
    .sync(FBHelper_sync)
  );
  assign io_in_fb_aw_ready = fb_io_in_aw_ready; // @[AXI4VGA.scala 130:15]
  assign io_in_fb_w_ready = fb_io_in_w_ready; // @[AXI4VGA.scala 131:14]
  assign io_in_fb_b_valid = fb_io_in_b_valid; // @[AXI4VGA.scala 132:14]
  assign io_in_fb_ar_ready = 1'h1; // @[AXI4VGA.scala 133:21]
  assign io_in_fb_r_valid = _T_2; // @[AXI4VGA.scala 136:20]
  assign io_in_ctrl_aw_ready = ctrl_io_in_aw_ready; // @[AXI4VGA.scala 126:14]
  assign io_in_ctrl_w_ready = ctrl_io_in_w_ready; // @[AXI4VGA.scala 126:14]
  assign io_in_ctrl_b_valid = ctrl_io_in_b_valid; // @[AXI4VGA.scala 126:14]
  assign io_in_ctrl_ar_ready = ctrl_io_in_ar_ready; // @[AXI4VGA.scala 126:14]
  assign io_in_ctrl_r_valid = ctrl_io_in_r_valid; // @[AXI4VGA.scala 126:14]
  assign io_in_ctrl_r_bits_data = ctrl_io_in_r_bits_data; // @[AXI4VGA.scala 126:14]
  assign io_vga_valid = hInRange & vInRange; // @[AXI4VGA.scala 148:16]
  assign ctrl_clock = clock;
  assign ctrl_reset = reset;
  assign ctrl_io_in_aw_valid = io_in_ctrl_aw_valid; // @[AXI4VGA.scala 126:14]
  assign ctrl_io_in_w_valid = io_in_ctrl_w_valid; // @[AXI4VGA.scala 126:14]
  assign ctrl_io_in_b_ready = io_in_ctrl_b_ready; // @[AXI4VGA.scala 126:14]
  assign ctrl_io_in_ar_valid = io_in_ctrl_ar_valid; // @[AXI4VGA.scala 126:14]
  assign ctrl_io_in_ar_bits_addr = io_in_ctrl_ar_bits_addr; // @[AXI4VGA.scala 126:14]
  assign ctrl_io_in_r_ready = io_in_ctrl_r_ready; // @[AXI4VGA.scala 126:14]
  assign fb_clock = clock;
  assign fb_reset = reset;
  assign fb_io_in_aw_valid = io_in_fb_aw_valid; // @[AXI4VGA.scala 130:15]
  assign fb_io_in_aw_bits_addr = io_in_fb_aw_bits_addr; // @[AXI4VGA.scala 130:15]
  assign fb_io_in_w_valid = io_in_fb_w_valid; // @[AXI4VGA.scala 131:14]
  assign fb_io_in_w_bits_data = io_in_fb_w_bits_data; // @[AXI4VGA.scala 131:14]
  assign fb_io_in_w_bits_strb = io_in_fb_w_bits_strb; // @[AXI4VGA.scala 131:14]
  assign fb_io_in_b_ready = io_in_fb_b_ready; // @[AXI4VGA.scala 132:14]
  assign fb_io_in_ar_valid = _T_34 & hCounterIs2; // @[AXI4VGA.scala 162:21]
  assign fb_io_in_ar_bits_addr = {{13'd0}, _T_33}; // @[AXI4VGA.scala 161:25]
  assign fb_io_in_r_ready = 1'h1; // @[AXI4VGA.scala 164:20]
  assign FBHelper_clk = clock; // @[AXI4VGA.scala 172:21]
  assign FBHelper_valid = io_vga_valid; // @[AXI4VGA.scala 173:23]
  assign FBHelper_pixel = hCounter[1] ? _GEN_14[63:32] : _GEN_14[31:0]; // @[AXI4VGA.scala 174:23]
  assign FBHelper_sync = ctrl_io_extra_sync; // @[AXI4VGA.scala 175:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  hCounter = _RAND_1[10:0];
  _RAND_2 = {1{`RANDOM}};
  vCounter = _RAND_2[9:0];
  _RAND_3 = {1{`RANDOM}};
  fbPixelAddrV0 = _RAND_3[16:0];
  _RAND_4 = {1{`RANDOM}};
  fbPixelAddrV1 = _RAND_4[16:0];
  _RAND_5 = {1{`RANDOM}};
  _T_34 = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  _T_38 = _RAND_6[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_2 <= 1'h0;
    end else begin
      _T_2 <= _GEN_1;
    end
    if (reset) begin
      hCounter <= 11'h0;
    end else if (hFinish) begin
      hCounter <= 11'h0;
    end else begin
      hCounter <= _T_5;
    end
    if (reset) begin
      vCounter <= 10'h0;
    end else if (hFinish) begin
      if (_T_6) begin
        vCounter <= 10'h0;
      end else begin
        vCounter <= _T_8;
      end
    end
    if (reset) begin
      fbPixelAddrV0 <= 17'h0;
    end else if (_T_22) begin
      if (_T_24) begin
        fbPixelAddrV0 <= 17'h0;
      end else begin
        fbPixelAddrV0 <= _T_26;
      end
    end
    if (reset) begin
      fbPixelAddrV1 <= 17'h0;
    end else if (_T_27) begin
      if (_T_29) begin
        fbPixelAddrV1 <= 17'h0;
      end else begin
        fbPixelAddrV1 <= _T_31;
      end
    end
    _T_34 <= _T_20 & hCounterIsOdd;
    if (reset) begin
      _T_38 <= 64'h0;
    end else if (_T_36) begin
      _T_38 <= fb_io_in_r_bits_data;
    end
  end
endmodule
module AXI4Flash(
  input         clock,
  input         reset,
  output        io_in_aw_ready,
  input         io_in_aw_valid,
  output        io_in_w_ready,
  input         io_in_w_valid,
  input         io_in_b_ready,
  output        io_in_b_valid,
  output        io_in_ar_ready,
  input         io_in_ar_valid,
  input  [31:0] io_in_ar_bits_addr,
  input         io_in_r_ready,
  output        io_in_r_valid,
  output [63:0] io_in_r_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  _T_30 = io_in_ar_ready & io_in_ar_valid; // @[Decoupled.scala 40:37]
  wire  _T_31 = io_in_r_ready & io_in_r_valid; // @[Decoupled.scala 40:37]
  reg  r_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_31 ? 1'h0 : r_busy; // @[StopWatch.scala 26:19]
  wire  _GEN_1 = _T_30 | _GEN_0; // @[StopWatch.scala 27:20]
  wire  _T_33 = ~r_busy; // @[AXI4Slave.scala 71:32]
  reg  ren; // @[AXI4Slave.scala 73:17]
  wire  _T_42 = _T_30 | r_busy; // @[AXI4Slave.scala 74:52]
  wire  _T_43 = ren & _T_42; // @[AXI4Slave.scala 74:35]
  reg  _T_45; // @[StopWatch.scala 24:20]
  wire  _GEN_2 = _T_31 ? 1'h0 : _T_45; // @[StopWatch.scala 26:19]
  wire  _GEN_3 = _T_43 | _GEN_2; // @[StopWatch.scala 27:20]
  wire  _T_46 = io_in_aw_ready & io_in_aw_valid; // @[Decoupled.scala 40:37]
  wire  _T_47 = io_in_b_ready & io_in_b_valid; // @[Decoupled.scala 40:37]
  reg  w_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_4 = _T_47 ? 1'h0 : w_busy; // @[StopWatch.scala 26:19]
  wire  _GEN_5 = _T_46 | _GEN_4; // @[StopWatch.scala 27:20]
  wire  _T_50 = io_in_w_ready & io_in_w_valid; // @[Decoupled.scala 40:37]
  reg  _T_53; // @[StopWatch.scala 24:20]
  wire  _GEN_6 = _T_47 ? 1'h0 : _T_53; // @[StopWatch.scala 26:19]
  wire  _GEN_7 = _T_50 | _GEN_6; // @[StopWatch.scala 27:20]
  wire  _T_88 = 13'h0 == io_in_ar_bits_addr[12:0]; // @[LookupTree.scala 24:34]
  wire  _T_89 = 13'h4 == io_in_ar_bits_addr[12:0]; // @[LookupTree.scala 24:34]
  wire  _T_90 = 13'h8 == io_in_ar_bits_addr[12:0]; // @[LookupTree.scala 24:34]
  wire [20:0] _T_91 = _T_88 ? 21'h10029b : 21'h0; // @[Mux.scala 27:72]
  wire [24:0] _T_92 = _T_89 ? 25'h1f29293 : 25'h0; // @[Mux.scala 27:72]
  wire [17:0] _T_93 = _T_90 ? 18'h28067 : 18'h0; // @[Mux.scala 27:72]
  wire [24:0] _GEN_9 = {{4'd0}, _T_91}; // @[Mux.scala 27:72]
  wire [24:0] _T_94 = _GEN_9 | _T_92; // @[Mux.scala 27:72]
  wire [24:0] _GEN_10 = {{7'd0}, _T_93}; // @[Mux.scala 27:72]
  wire [24:0] _T_95 = _T_94 | _GEN_10; // @[Mux.scala 27:72]
  wire [63:0] rdata = {{39'd0}, _T_95}; // @[AXI4Flash.scala 37:19 RegMap.scala 30:11]
  reg [63:0] _T_99; // @[AXI4Flash.scala 41:38]
  reg [63:0] _T_100; // @[Reg.scala 15:16]
  assign io_in_aw_ready = ~w_busy; // @[AXI4Slave.scala 94:15]
  assign io_in_w_ready = io_in_aw_valid | w_busy; // @[AXI4Slave.scala 95:15]
  assign io_in_b_valid = _T_53; // @[AXI4Slave.scala 97:14]
  assign io_in_ar_ready = io_in_r_ready | _T_33; // @[AXI4Slave.scala 71:15]
  assign io_in_r_valid = _T_45; // @[AXI4Slave.scala 74:14]
  assign io_in_r_bits_data = _T_100; // @[AXI4Flash.scala 41:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ren = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _T_45 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_53 = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  _T_99 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  _T_100 = _RAND_6[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      r_busy <= 1'h0;
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin
      ren <= 1'h0;
    end else begin
      ren <= _T_30;
    end
    if (reset) begin
      _T_45 <= 1'h0;
    end else begin
      _T_45 <= _GEN_3;
    end
    if (reset) begin
      w_busy <= 1'h0;
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin
      _T_53 <= 1'h0;
    end else begin
      _T_53 <= _GEN_7;
    end
    _T_99 <= {rdata[31:0],rdata[31:0]};
    if (ren) begin
      _T_100 <= _T_99;
    end
  end
endmodule
module AXI4DummySD(
  input         clock,
  input         reset,
  output        io_in_aw_ready,
  input         io_in_aw_valid,
  input  [31:0] io_in_aw_bits_addr,
  output        io_in_w_ready,
  input         io_in_w_valid,
  input  [63:0] io_in_w_bits_data,
  input  [7:0]  io_in_w_bits_strb,
  input         io_in_b_ready,
  output        io_in_b_valid,
  output        io_in_ar_ready,
  input         io_in_ar_valid,
  input  [31:0] io_in_ar_bits_addr,
  input         io_in_r_ready,
  output        io_in_r_valid,
  output [63:0] io_in_r_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  wire  sdHelper_clk; // @[AXI4DummySD.scala 114:24]
  wire  sdHelper_ren; // @[AXI4DummySD.scala 114:24]
  wire [31:0] sdHelper_data; // @[AXI4DummySD.scala 114:24]
  wire  sdHelper_setAddr; // @[AXI4DummySD.scala 114:24]
  wire [31:0] sdHelper_addr; // @[AXI4DummySD.scala 114:24]
  wire  _T_30 = io_in_ar_ready & io_in_ar_valid; // @[Decoupled.scala 40:37]
  wire  _T_31 = io_in_r_ready & io_in_r_valid; // @[Decoupled.scala 40:37]
  reg  r_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_31 ? 1'h0 : r_busy; // @[StopWatch.scala 26:19]
  wire  _GEN_1 = _T_30 | _GEN_0; // @[StopWatch.scala 27:20]
  wire  _T_33 = ~r_busy; // @[AXI4Slave.scala 71:32]
  reg  ren; // @[AXI4Slave.scala 73:17]
  wire  _T_42 = _T_30 | r_busy; // @[AXI4Slave.scala 74:52]
  wire  _T_43 = ren & _T_42; // @[AXI4Slave.scala 74:35]
  reg  _T_45; // @[StopWatch.scala 24:20]
  wire  _GEN_2 = _T_31 ? 1'h0 : _T_45; // @[StopWatch.scala 26:19]
  wire  _GEN_3 = _T_43 | _GEN_2; // @[StopWatch.scala 27:20]
  wire  _T_46 = io_in_aw_ready & io_in_aw_valid; // @[Decoupled.scala 40:37]
  wire  _T_47 = io_in_b_ready & io_in_b_valid; // @[Decoupled.scala 40:37]
  reg  w_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_4 = _T_47 ? 1'h0 : w_busy; // @[StopWatch.scala 26:19]
  wire  _GEN_5 = _T_46 | _GEN_4; // @[StopWatch.scala 27:20]
  wire  _T_50 = io_in_w_ready & io_in_w_valid; // @[Decoupled.scala 40:37]
  reg  _T_53; // @[StopWatch.scala 24:20]
  wire  _GEN_6 = _T_47 ? 1'h0 : _T_53; // @[StopWatch.scala 26:19]
  wire  _GEN_7 = _T_50 | _GEN_6; // @[StopWatch.scala 27:20]
  reg [31:0] regs_0; // @[AXI4DummySD.scala 72:43]
  reg [31:0] regs_1; // @[AXI4DummySD.scala 72:43]
  reg [31:0] regs_4; // @[AXI4DummySD.scala 72:43]
  reg [31:0] regs_5; // @[AXI4DummySD.scala 72:43]
  reg [31:0] regs_6; // @[AXI4DummySD.scala 72:43]
  reg [31:0] regs_7; // @[AXI4DummySD.scala 72:43]
  reg [31:0] regs_8; // @[AXI4DummySD.scala 72:43]
  reg [31:0] regs_15; // @[AXI4DummySD.scala 72:43]
  reg [31:0] regs_20; // @[AXI4DummySD.scala 72:43]
  wire  _T_55 = io_in_ar_bits_addr[12:0] == 13'h40; // @[AXI4DummySD.scala 116:40]
  wire [3:0] strb = io_in_aw_bits_addr[2] ? io_in_w_bits_strb[7:4] : io_in_w_bits_strb[3:0]; // @[AXI4DummySD.scala 138:22]
  wire [7:0] _T_69 = strb[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_71 = strb[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_73 = strb[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_75 = strb[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_78 = {_T_75,_T_73,_T_71,_T_69}; // @[Cat.scala 29:58]
  wire  _T_79 = 13'h0 == io_in_ar_bits_addr[12:0]; // @[LookupTree.scala 24:34]
  wire  _T_80 = 13'h38 == io_in_ar_bits_addr[12:0]; // @[LookupTree.scala 24:34]
  wire  _T_81 = 13'h18 == io_in_ar_bits_addr[12:0]; // @[LookupTree.scala 24:34]
  wire  _T_82 = 13'h34 == io_in_ar_bits_addr[12:0]; // @[LookupTree.scala 24:34]
  wire  _T_83 = 13'h14 == io_in_ar_bits_addr[12:0]; // @[LookupTree.scala 24:34]
  wire  _T_84 = 13'h1c == io_in_ar_bits_addr[12:0]; // @[LookupTree.scala 24:34]
  wire  _T_85 = 13'h20 == io_in_ar_bits_addr[12:0]; // @[LookupTree.scala 24:34]
  wire  _T_86 = 13'h40 == io_in_ar_bits_addr[12:0]; // @[LookupTree.scala 24:34]
  wire  _T_87 = 13'h50 == io_in_ar_bits_addr[12:0]; // @[LookupTree.scala 24:34]
  wire  _T_88 = 13'h10 == io_in_ar_bits_addr[12:0]; // @[LookupTree.scala 24:34]
  wire  _T_89 = 13'h4 == io_in_ar_bits_addr[12:0]; // @[LookupTree.scala 24:34]
  wire [31:0] _T_90 = _T_79 ? regs_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_91 = _T_80 ? regs_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_92 = _T_81 ? regs_6 : 32'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_93 = _T_82 ? 8'h80 : 8'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_94 = _T_83 ? regs_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_95 = _T_84 ? regs_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_96 = _T_85 ? regs_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_97 = _T_86 ? sdHelper_data : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_98 = _T_87 ? regs_20 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_99 = _T_88 ? regs_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_100 = _T_89 ? regs_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_101 = _T_90 | _T_91; // @[Mux.scala 27:72]
  wire [31:0] _T_102 = _T_101 | _T_92; // @[Mux.scala 27:72]
  wire [31:0] _GEN_40 = {{24'd0}, _T_93}; // @[Mux.scala 27:72]
  wire [31:0] _T_103 = _T_102 | _GEN_40; // @[Mux.scala 27:72]
  wire [31:0] _T_104 = _T_103 | _T_94; // @[Mux.scala 27:72]
  wire [31:0] _T_105 = _T_104 | _T_95; // @[Mux.scala 27:72]
  wire [31:0] _T_106 = _T_105 | _T_96; // @[Mux.scala 27:72]
  wire [31:0] _T_107 = _T_106 | _T_97; // @[Mux.scala 27:72]
  wire [31:0] _T_108 = _T_107 | _T_98; // @[Mux.scala 27:72]
  wire [31:0] _T_109 = _T_108 | _T_99; // @[Mux.scala 27:72]
  wire [31:0] _T_110 = _T_109 | _T_100; // @[Mux.scala 27:72]
  wire  _T_112 = io_in_aw_bits_addr[12:0] == 13'h0; // @[RegMap.scala 32:41]
  wire  _T_113 = _T_50 & _T_112; // @[RegMap.scala 32:32]
  wire [63:0] _GEN_41 = {{32'd0}, _T_78}; // @[BitUtils.scala 32:13]
  wire [63:0] _T_114 = io_in_w_bits_data & _GEN_41; // @[BitUtils.scala 32:13]
  wire [31:0] _T_115 = ~_T_78; // @[BitUtils.scala 32:38]
  wire [31:0] _T_116 = regs_0 & _T_115; // @[BitUtils.scala 32:36]
  wire [63:0] _GEN_42 = {{32'd0}, _T_116}; // @[BitUtils.scala 32:25]
  wire [63:0] _T_117 = _T_114 | _GEN_42; // @[BitUtils.scala 32:25]
  wire  _T_119 = 6'h1 == _T_117[5:0]; // @[Conditional.scala 37:30]
  wire  _T_120 = 6'h2 == _T_117[5:0]; // @[Conditional.scala 37:30]
  wire  _T_121 = 6'h9 == _T_117[5:0]; // @[Conditional.scala 37:30]
  wire  _T_127 = 6'hd == _T_117[5:0]; // @[Conditional.scala 37:30]
  wire  _T_128 = 6'h12 == _T_117[5:0]; // @[Conditional.scala 37:30]
  wire  _GEN_13 = _T_127 ? 1'h0 : _T_128; // @[Conditional.scala 39:67]
  wire  _GEN_18 = _T_121 ? 1'h0 : _GEN_13; // @[Conditional.scala 39:67]
  wire  _GEN_23 = _T_120 ? 1'h0 : _GEN_18; // @[Conditional.scala 39:67]
  wire  _GEN_28 = _T_119 ? 1'h0 : _GEN_23; // @[Conditional.scala 40:58]
  wire [63:0] _GEN_34 = _T_113 ? _T_117 : {{32'd0}, regs_0}; // @[RegMap.scala 32:48]
  wire  _T_129 = io_in_aw_bits_addr[12:0] == 13'h38; // @[RegMap.scala 32:41]
  wire  _T_130 = _T_50 & _T_129; // @[RegMap.scala 32:32]
  wire [31:0] _T_133 = regs_15 & _T_115; // @[BitUtils.scala 32:36]
  wire [63:0] _GEN_44 = {{32'd0}, _T_133}; // @[BitUtils.scala 32:25]
  wire [63:0] _T_134 = _T_114 | _GEN_44; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_35 = _T_130 ? _T_134 : {{32'd0}, regs_15}; // @[RegMap.scala 32:48]
  wire  _T_135 = io_in_aw_bits_addr[12:0] == 13'h20; // @[RegMap.scala 32:41]
  wire  _T_136 = _T_50 & _T_135; // @[RegMap.scala 32:32]
  wire [31:0] _T_139 = regs_8 & _T_115; // @[BitUtils.scala 32:36]
  wire [63:0] _GEN_46 = {{32'd0}, _T_139}; // @[BitUtils.scala 32:25]
  wire [63:0] _T_140 = _T_114 | _GEN_46; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_36 = _T_136 ? _T_140 : {{32'd0}, regs_8}; // @[RegMap.scala 32:48]
  wire  _T_141 = io_in_aw_bits_addr[12:0] == 13'h50; // @[RegMap.scala 32:41]
  wire  _T_142 = _T_50 & _T_141; // @[RegMap.scala 32:32]
  wire [31:0] _T_145 = regs_20 & _T_115; // @[BitUtils.scala 32:36]
  wire [63:0] _GEN_48 = {{32'd0}, _T_145}; // @[BitUtils.scala 32:25]
  wire [63:0] _T_146 = _T_114 | _GEN_48; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_37 = _T_142 ? _T_146 : {{32'd0}, regs_20}; // @[RegMap.scala 32:48]
  wire  _T_147 = io_in_aw_bits_addr[12:0] == 13'h4; // @[RegMap.scala 32:41]
  wire  _T_148 = _T_50 & _T_147; // @[RegMap.scala 32:32]
  wire [31:0] _T_151 = regs_1 & _T_115; // @[BitUtils.scala 32:36]
  wire [63:0] _GEN_50 = {{32'd0}, _T_151}; // @[BitUtils.scala 32:25]
  wire [63:0] _T_152 = _T_114 | _GEN_50; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_38 = _T_148 ? _T_152 : {{32'd0}, regs_1}; // @[RegMap.scala 32:48]
  wire [63:0] rdata = {{32'd0}, _T_110}; // @[AXI4DummySD.scala 139:19 RegMap.scala 30:11]
  reg [63:0] _T_155; // @[AXI4DummySD.scala 144:44]
  reg [63:0] _T_156; // @[Reg.scala 15:16]
  SDHelper sdHelper ( // @[AXI4DummySD.scala 114:24]
    .clk(sdHelper_clk),
    .ren(sdHelper_ren),
    .data(sdHelper_data),
    .setAddr(sdHelper_setAddr),
    .addr(sdHelper_addr)
  );
  assign io_in_aw_ready = ~w_busy; // @[AXI4Slave.scala 94:15]
  assign io_in_w_ready = io_in_aw_valid | w_busy; // @[AXI4Slave.scala 95:15]
  assign io_in_b_valid = _T_53; // @[AXI4Slave.scala 97:14]
  assign io_in_ar_ready = io_in_r_ready | _T_33; // @[AXI4Slave.scala 71:15]
  assign io_in_r_valid = _T_45; // @[AXI4Slave.scala 74:14]
  assign io_in_r_bits_data = _T_156; // @[AXI4DummySD.scala 143:18]
  assign sdHelper_clk = clock; // @[AXI4DummySD.scala 115:19]
  assign sdHelper_ren = _T_55 & _T_30; // @[AXI4DummySD.scala 116:19]
  assign sdHelper_setAddr = _T_113 & _GEN_28; // @[AXI4DummySD.scala 117:23]
  assign sdHelper_addr = regs_1; // @[AXI4DummySD.scala 118:20]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ren = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _T_45 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_53 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  regs_0 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  regs_1 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  regs_4 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  regs_5 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  regs_6 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  regs_7 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  regs_8 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  regs_15 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  regs_20 = _RAND_13[31:0];
  _RAND_14 = {2{`RANDOM}};
  _T_155 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  _T_156 = _RAND_15[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      r_busy <= 1'h0;
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin
      ren <= 1'h0;
    end else begin
      ren <= _T_30;
    end
    if (reset) begin
      _T_45 <= 1'h0;
    end else begin
      _T_45 <= _GEN_3;
    end
    if (reset) begin
      w_busy <= 1'h0;
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin
      _T_53 <= 1'h0;
    end else begin
      _T_53 <= _GEN_7;
    end
    if (reset) begin
      regs_0 <= 32'h0;
    end else begin
      regs_0 <= _GEN_34[31:0];
    end
    if (reset) begin
      regs_1 <= 32'h0;
    end else begin
      regs_1 <= _GEN_38[31:0];
    end
    if (reset) begin
      regs_4 <= 32'h0;
    end else if (_T_113) begin
      if (_T_119) begin
        regs_4 <= 32'h80ff8000;
      end else if (_T_120) begin
        regs_4 <= 32'h1;
      end else if (_T_121) begin
        regs_4 <= 32'h92404001;
      end else if (_T_127) begin
        regs_4 <= 32'h0;
      end
    end
    if (reset) begin
      regs_5 <= 32'h0;
    end else if (_T_113) begin
      if (!(_T_119)) begin
        if (_T_120) begin
          regs_5 <= 32'h0;
        end else if (_T_121) begin
          regs_5 <= 32'hd24b97e3;
        end else if (_T_127) begin
          regs_5 <= 32'h0;
        end
      end
    end
    if (reset) begin
      regs_6 <= 32'h0;
    end else if (_T_113) begin
      if (!(_T_119)) begin
        if (_T_120) begin
          regs_6 <= 32'h0;
        end else if (_T_121) begin
          regs_6 <= 32'hf5f803f;
        end else if (_T_127) begin
          regs_6 <= 32'h0;
        end
      end
    end
    if (reset) begin
      regs_7 <= 32'h0;
    end else if (_T_113) begin
      if (!(_T_119)) begin
        if (_T_120) begin
          regs_7 <= 32'h15000000;
        end else if (_T_121) begin
          regs_7 <= 32'h8c26012a;
        end else if (_T_127) begin
          regs_7 <= 32'h0;
        end
      end
    end
    if (reset) begin
      regs_8 <= 32'h0;
    end else begin
      regs_8 <= _GEN_36[31:0];
    end
    if (reset) begin
      regs_15 <= 32'h0;
    end else begin
      regs_15 <= _GEN_35[31:0];
    end
    if (reset) begin
      regs_20 <= 32'h0;
    end else begin
      regs_20 <= _GEN_37[31:0];
    end
    _T_155 <= {rdata[31:0],rdata[31:0]};
    if (ren) begin
      _T_156 <= _T_155;
    end
  end
endmodule
module AXI4DiffTestCtrl(
  input         clock,
  input         reset,
  output        io_in_aw_ready,
  input         io_in_aw_valid,
  input  [31:0] io_in_aw_bits_addr,
  output        io_in_w_ready,
  input         io_in_w_valid,
  input  [63:0] io_in_w_bits_data,
  input  [7:0]  io_in_w_bits_strb,
  input         io_in_b_ready,
  output        io_in_b_valid,
  output        io_in_ar_ready,
  input         io_in_ar_valid,
  input         io_in_r_ready,
  output        io_in_r_valid,
  output [63:0] io_in_r_bits_data,
  output        io_extra_enable
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] _T_9 = io_in_w_bits_strb[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_11 = io_in_w_bits_strb[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_13 = io_in_w_bits_strb[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_15 = io_in_w_bits_strb[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_17 = io_in_w_bits_strb[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_19 = io_in_w_bits_strb[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_21 = io_in_w_bits_strb[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_23 = io_in_w_bits_strb[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] fullMask = {_T_23,_T_21,_T_19,_T_17,_T_15,_T_13,_T_11,_T_9}; // @[Cat.scala 29:58]
  wire  _T_30 = io_in_ar_ready & io_in_ar_valid; // @[Decoupled.scala 40:37]
  wire  _T_31 = io_in_r_ready & io_in_r_valid; // @[Decoupled.scala 40:37]
  reg  r_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_31 ? 1'h0 : r_busy; // @[StopWatch.scala 26:19]
  wire  _GEN_1 = _T_30 | _GEN_0; // @[StopWatch.scala 27:20]
  wire  _T_33 = ~r_busy; // @[AXI4Slave.scala 71:32]
  reg  ren; // @[AXI4Slave.scala 73:17]
  wire  _T_42 = _T_30 | r_busy; // @[AXI4Slave.scala 74:52]
  wire  _T_43 = ren & _T_42; // @[AXI4Slave.scala 74:35]
  reg  _T_45; // @[StopWatch.scala 24:20]
  wire  _GEN_2 = _T_31 ? 1'h0 : _T_45; // @[StopWatch.scala 26:19]
  wire  _GEN_3 = _T_43 | _GEN_2; // @[StopWatch.scala 27:20]
  wire  _T_46 = io_in_aw_ready & io_in_aw_valid; // @[Decoupled.scala 40:37]
  wire  _T_47 = io_in_b_ready & io_in_b_valid; // @[Decoupled.scala 40:37]
  reg  w_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_4 = _T_47 ? 1'h0 : w_busy; // @[StopWatch.scala 26:19]
  wire  _GEN_5 = _T_46 | _GEN_4; // @[StopWatch.scala 27:20]
  wire  _T_50 = io_in_w_ready & io_in_w_valid; // @[Decoupled.scala 40:37]
  reg  _T_53; // @[StopWatch.scala 24:20]
  wire  _GEN_6 = _T_47 ? 1'h0 : _T_53; // @[StopWatch.scala 26:19]
  wire  _GEN_7 = _T_50 | _GEN_6; // @[StopWatch.scala 27:20]
  reg  enable; // @[DiffTest.scala 31:23]
  wire  _T_89 = io_in_aw_bits_addr[3:0] == 4'h0; // @[RegMap.scala 32:41]
  wire  _T_90 = _T_50 & _T_89; // @[RegMap.scala 32:32]
  wire [63:0] _T_91 = io_in_w_bits_data & fullMask; // @[BitUtils.scala 32:13]
  wire [63:0] _T_92 = ~fullMask; // @[BitUtils.scala 32:38]
  wire [63:0] _GEN_9 = {{63'd0}, enable}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_93 = _GEN_9 & _T_92; // @[BitUtils.scala 32:36]
  wire [63:0] _T_94 = _T_91 | _T_93; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_8 = _T_90 ? _T_94 : {{63'd0}, enable}; // @[RegMap.scala 32:48]
  assign io_in_aw_ready = ~w_busy; // @[AXI4Slave.scala 94:15]
  assign io_in_w_ready = io_in_aw_valid | w_busy; // @[AXI4Slave.scala 95:15]
  assign io_in_b_valid = _T_53; // @[AXI4Slave.scala 97:14]
  assign io_in_ar_ready = io_in_r_ready | _T_33; // @[AXI4Slave.scala 71:15]
  assign io_in_r_valid = _T_45; // @[AXI4Slave.scala 74:14]
  assign io_in_r_bits_data = {{63'd0}, enable}; // @[RegMap.scala 30:11]
  assign io_extra_enable = enable; // @[DiffTest.scala 41:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ren = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _T_45 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_53 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  enable = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      r_busy <= 1'h0;
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin
      ren <= 1'h0;
    end else begin
      ren <= _T_30;
    end
    if (reset) begin
      _T_45 <= 1'h0;
    end else begin
      _T_45 <= _GEN_3;
    end
    if (reset) begin
      w_busy <= 1'h0;
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin
      _T_53 <= 1'h0;
    end else begin
      _T_53 <= _GEN_7;
    end
    if (reset) begin
      enable <= 1'h0;
    end else begin
      enable <= _GEN_8[0];
    end
  end
endmodule
module AXI4DMA(
  input         clock,
  input         reset,
  output        io_in_aw_ready,
  input         io_in_aw_valid,
  input  [31:0] io_in_aw_bits_addr,
  output        io_in_w_ready,
  input         io_in_w_valid,
  input  [63:0] io_in_w_bits_data,
  input  [7:0]  io_in_w_bits_strb,
  input         io_in_b_ready,
  output        io_in_b_valid,
  output        io_in_ar_ready,
  input         io_in_ar_valid,
  input  [31:0] io_in_ar_bits_addr,
  input         io_in_r_ready,
  output        io_in_r_valid,
  output [63:0] io_in_r_bits_data,
  input         io_extra_dma_aw_ready,
  output        io_extra_dma_aw_valid,
  output [31:0] io_extra_dma_aw_bits_addr,
  output [7:0]  io_extra_dma_aw_bits_len,
  output [2:0]  io_extra_dma_aw_bits_size,
  input         io_extra_dma_w_ready,
  output        io_extra_dma_w_valid,
  output [63:0] io_extra_dma_w_bits_data,
  output [7:0]  io_extra_dma_w_bits_strb,
  output        io_extra_dma_w_bits_last,
  output        io_extra_dma_b_ready,
  input         io_extra_dma_b_valid,
  input         io_extra_dma_ar_ready,
  output        io_extra_dma_ar_valid,
  output [31:0] io_extra_dma_ar_bits_addr,
  output [7:0]  io_extra_dma_ar_bits_len,
  output [2:0]  io_extra_dma_ar_bits_size,
  output        io_extra_dma_r_ready,
  input         io_extra_dma_r_valid,
  input  [63:0] io_extra_dma_r_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire  _T_30 = io_in_ar_ready & io_in_ar_valid; // @[Decoupled.scala 40:37]
  wire  _T_31 = io_in_r_ready & io_in_r_valid; // @[Decoupled.scala 40:37]
  reg  r_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_31 ? 1'h0 : r_busy; // @[StopWatch.scala 26:19]
  wire  _GEN_1 = _T_30 | _GEN_0; // @[StopWatch.scala 27:20]
  wire  _T_33 = ~r_busy; // @[AXI4Slave.scala 71:32]
  reg  ren; // @[AXI4Slave.scala 73:17]
  wire  _T_42 = _T_30 | r_busy; // @[AXI4Slave.scala 74:52]
  wire  _T_43 = ren & _T_42; // @[AXI4Slave.scala 74:35]
  reg  _T_45; // @[StopWatch.scala 24:20]
  wire  _GEN_2 = _T_31 ? 1'h0 : _T_45; // @[StopWatch.scala 26:19]
  wire  _GEN_3 = _T_43 | _GEN_2; // @[StopWatch.scala 27:20]
  wire  _T_46 = io_in_aw_ready & io_in_aw_valid; // @[Decoupled.scala 40:37]
  wire  _T_47 = io_in_b_ready & io_in_b_valid; // @[Decoupled.scala 40:37]
  reg  w_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_4 = _T_47 ? 1'h0 : w_busy; // @[StopWatch.scala 26:19]
  wire  _GEN_5 = _T_46 | _GEN_4; // @[StopWatch.scala 27:20]
  wire  _T_50 = io_in_w_ready & io_in_w_valid; // @[Decoupled.scala 40:37]
  reg  _T_53; // @[StopWatch.scala 24:20]
  wire  _GEN_6 = _T_47 ? 1'h0 : _T_53; // @[StopWatch.scala 26:19]
  wire  _GEN_7 = _T_50 | _GEN_6; // @[StopWatch.scala 27:20]
  reg [31:0] dest; // @[AXI4DMA.scala 34:17]
  reg [31:0] src; // @[AXI4DMA.scala 35:16]
  reg [31:0] len; // @[AXI4DMA.scala 36:20]
  reg [31:0] data; // @[AXI4DMA.scala 39:17]
  reg [2:0] state; // @[AXI4DMA.scala 42:22]
  wire  _T_54 = state == 3'h0; // @[AXI4DMA.scala 52:15]
  wire  _T_55 = len != 32'h0; // @[AXI4DMA.scala 52:33]
  wire  _T_56 = _T_54 & _T_55; // @[AXI4DMA.scala 52:26]
  wire  _T_57 = state == 3'h1; // @[AXI4DMA.scala 53:15]
  wire  _T_58 = io_extra_dma_ar_ready & io_extra_dma_ar_valid; // @[Decoupled.scala 40:37]
  wire  _T_59 = _T_57 & _T_58; // @[AXI4DMA.scala 53:30]
  wire  _T_60 = state == 3'h2; // @[AXI4DMA.scala 54:15]
  wire  _T_61 = io_extra_dma_r_ready & io_extra_dma_r_valid; // @[Decoupled.scala 40:37]
  wire  _T_62 = _T_60 & _T_61; // @[AXI4DMA.scala 54:36]
  wire  _T_68 = io_extra_dma_aw_ready & io_extra_dma_aw_valid; // @[Decoupled.scala 40:37]
  reg  awAck; // @[StopWatch.scala 24:20]
  wire  _GEN_14 = _T_68 | awAck; // @[StopWatch.scala 30:20]
  wire  _T_72 = io_extra_dma_w_ready & io_extra_dma_w_valid; // @[Decoupled.scala 40:37]
  wire  _T_73 = _T_68 & _T_72; // @[AXI4DMA.scala 63:27]
  wire  _T_74 = _T_73 & io_extra_dma_w_bits_last; // @[AXI4DMA.scala 63:43]
  reg  wAck; // @[StopWatch.scala 24:20]
  wire  _T_75 = awAck & wAck; // @[AXI4DMA.scala 63:63]
  wire  wSend = _T_74 | _T_75; // @[AXI4DMA.scala 63:53]
  wire  _T_70 = _T_72 & io_extra_dma_w_bits_last; // @[AXI4DMA.scala 62:41]
  wire  _GEN_16 = _T_70 | wAck; // @[StopWatch.scala 30:20]
  wire  _T_77 = state == 3'h3; // @[AXI4DMA.scala 65:15]
  wire  _T_78 = _T_77 & wSend; // @[AXI4DMA.scala 65:31]
  wire  _T_79 = state == 3'h4; // @[AXI4DMA.scala 66:15]
  wire  _T_80 = io_extra_dma_b_ready & io_extra_dma_b_valid; // @[Decoupled.scala 40:37]
  wire  _T_81 = _T_79 & _T_80; // @[AXI4DMA.scala 66:37]
  wire [31:0] _T_83 = len - 32'h4; // @[AXI4DMA.scala 67:16]
  wire [31:0] _T_85 = dest + 32'h4; // @[AXI4DMA.scala 68:18]
  wire [31:0] _T_87 = src + 32'h4; // @[AXI4DMA.scala 69:16]
  wire  _T_88 = len <= 32'h4; // @[AXI4DMA.scala 70:22]
  wire [31:0] _GEN_19 = _T_81 ? _T_83 : len; // @[AXI4DMA.scala 66:54]
  wire [31:0] _GEN_20 = _T_81 ? _T_85 : dest; // @[AXI4DMA.scala 66:54]
  wire [31:0] _GEN_21 = _T_81 ? _T_87 : src; // @[AXI4DMA.scala 66:54]
  wire  _T_93 = ~awAck; // @[AXI4DMA.scala 88:46]
  wire  _T_96 = ~wAck; // @[AXI4DMA.scala 89:45]
  wire [2:0] _GEN_26 = {{2'd0}, dest[2]}; // @[AXI4DMA.scala 91:68]
  wire [3:0] _T_101 = _GEN_26 * 3'h4; // @[AXI4DMA.scala 91:68]
  wire [18:0] _T_102 = 19'hf << _T_101; // @[AXI4DMA.scala 91:41]
  wire [7:0] _T_108 = io_in_w_bits_strb >> io_in_aw_bits_addr[2:0]; // @[AXI4DMA.scala 102:72]
  wire [7:0] _T_118 = _T_108[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_120 = _T_108[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_122 = _T_108[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_124 = _T_108[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_126 = _T_108[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_128 = _T_108[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_130 = _T_108[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_132 = _T_108[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_139 = {_T_132,_T_130,_T_128,_T_126,_T_124,_T_122,_T_120,_T_118}; // @[Cat.scala 29:58]
  wire  _T_140 = 4'h0 == io_in_ar_bits_addr[3:0]; // @[LookupTree.scala 24:34]
  wire  _T_141 = 4'h4 == io_in_ar_bits_addr[3:0]; // @[LookupTree.scala 24:34]
  wire  _T_142 = 4'h8 == io_in_ar_bits_addr[3:0]; // @[LookupTree.scala 24:34]
  wire [31:0] _T_143 = _T_140 ? dest : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_144 = _T_141 ? src : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_145 = _T_142 ? len : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_146 = _T_143 | _T_144; // @[Mux.scala 27:72]
  wire [31:0] _T_147 = _T_146 | _T_145; // @[Mux.scala 27:72]
  wire  _T_149 = io_in_aw_bits_addr[3:0] == 4'h0; // @[RegMap.scala 32:41]
  wire  _T_150 = _T_50 & _T_149; // @[RegMap.scala 32:32]
  wire [63:0] _T_151 = io_in_w_bits_data & _T_139; // @[BitUtils.scala 32:13]
  wire [63:0] _T_152 = ~_T_139; // @[BitUtils.scala 32:38]
  wire [63:0] _GEN_27 = {{32'd0}, dest}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_153 = _GEN_27 & _T_152; // @[BitUtils.scala 32:36]
  wire [63:0] _T_154 = _T_151 | _T_153; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_23 = _T_150 ? _T_154 : {{32'd0}, _GEN_20}; // @[RegMap.scala 32:48]
  wire  _T_155 = io_in_aw_bits_addr[3:0] == 4'h4; // @[RegMap.scala 32:41]
  wire  _T_156 = _T_50 & _T_155; // @[RegMap.scala 32:32]
  wire [63:0] _GEN_28 = {{32'd0}, src}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_159 = _GEN_28 & _T_152; // @[BitUtils.scala 32:36]
  wire [63:0] _T_160 = _T_151 | _T_159; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_24 = _T_156 ? _T_160 : {{32'd0}, _GEN_21}; // @[RegMap.scala 32:48]
  wire  _T_161 = io_in_aw_bits_addr[3:0] == 4'h8; // @[RegMap.scala 32:41]
  wire  _T_162 = _T_50 & _T_161; // @[RegMap.scala 32:32]
  wire [63:0] _GEN_29 = {{32'd0}, len}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_165 = _GEN_29 & _T_152; // @[BitUtils.scala 32:36]
  wire [63:0] _T_166 = _T_151 | _T_165; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_25 = _T_162 ? _T_166 : {{32'd0}, _GEN_19}; // @[RegMap.scala 32:48]
  assign io_in_aw_ready = ~w_busy; // @[AXI4Slave.scala 94:15]
  assign io_in_w_ready = io_in_aw_valid | w_busy; // @[AXI4Slave.scala 95:15]
  assign io_in_b_valid = _T_53; // @[AXI4Slave.scala 97:14]
  assign io_in_ar_ready = io_in_r_ready | _T_33; // @[AXI4Slave.scala 71:15]
  assign io_in_r_valid = _T_45; // @[AXI4Slave.scala 74:14]
  assign io_in_r_bits_data = {{32'd0}, _T_147}; // @[RegMap.scala 30:11]
  assign io_extra_dma_aw_valid = _T_77 & _T_93; // @[AXI4DMA.scala 88:16]
  assign io_extra_dma_aw_bits_addr = dest; // @[AXI4DMA.scala 86:15 AXI4DMA.scala 87:20]
  assign io_extra_dma_aw_bits_len = io_extra_dma_ar_bits_len; // @[AXI4DMA.scala 86:15]
  assign io_extra_dma_aw_bits_size = io_extra_dma_ar_bits_size; // @[AXI4DMA.scala 86:15]
  assign io_extra_dma_w_valid = _T_77 & _T_96; // @[AXI4DMA.scala 89:15]
  assign io_extra_dma_w_bits_data = {data,data}; // @[AXI4DMA.scala 90:19]
  assign io_extra_dma_w_bits_strb = _T_102[7:0]; // @[AXI4DMA.scala 91:19]
  assign io_extra_dma_w_bits_last = 1'h1; // @[AXI4DMA.scala 92:19]
  assign io_extra_dma_b_ready = state == 3'h4; // @[AXI4DMA.scala 93:15]
  assign io_extra_dma_ar_valid = state == 3'h1; // @[AXI4DMA.scala 83:16]
  assign io_extra_dma_ar_bits_addr = src; // @[AXI4DMA.scala 82:20]
  assign io_extra_dma_ar_bits_len = 8'h0; // @[AXI4DMA.scala 81:19]
  assign io_extra_dma_ar_bits_size = 3'h2; // @[AXI4DMA.scala 75:20]
  assign io_extra_dma_r_ready = state == 3'h2; // @[AXI4DMA.scala 84:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ren = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _T_45 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_53 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  dest = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  src = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  len = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  data = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  state = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  awAck = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  wAck = _RAND_11[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      r_busy <= 1'h0;
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin
      ren <= 1'h0;
    end else begin
      ren <= _T_30;
    end
    if (reset) begin
      _T_45 <= 1'h0;
    end else begin
      _T_45 <= _GEN_3;
    end
    if (reset) begin
      w_busy <= 1'h0;
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin
      _T_53 <= 1'h0;
    end else begin
      _T_53 <= _GEN_7;
    end
    dest <= _GEN_23[31:0];
    src <= _GEN_24[31:0];
    if (reset) begin
      len <= 32'h0;
    end else begin
      len <= _GEN_25[31:0];
    end
    if (_T_62) begin
      if (src[2]) begin
        data <= io_extra_dma_r_bits_data[63:32];
      end else begin
        data <= io_extra_dma_r_bits_data[31:0];
      end
    end
    if (reset) begin
      state <= 3'h0;
    end else if (_T_81) begin
      if (_T_88) begin
        state <= 3'h0;
      end else begin
        state <= 3'h1;
      end
    end else if (_T_78) begin
      state <= 3'h4;
    end else if (_T_62) begin
      state <= 3'h3;
    end else if (_T_59) begin
      state <= 3'h2;
    end else if (_T_56) begin
      state <= 3'h1;
    end
    if (reset) begin
      awAck <= 1'h0;
    end else if (wSend) begin
      awAck <= 1'h0;
    end else begin
      awAck <= _GEN_14;
    end
    if (reset) begin
      wAck <= 1'h0;
    end else if (wSend) begin
      wAck <= 1'h0;
    end else begin
      wAck <= _GEN_16;
    end
  end
endmodule
module SimMMIO(
  input         clock,
  input         reset,
  output        io_rw_req_ready,
  input         io_rw_req_valid,
  input  [31:0] io_rw_req_bits_addr,
  input  [2:0]  io_rw_req_bits_size,
  input  [3:0]  io_rw_req_bits_cmd,
  input  [7:0]  io_rw_req_bits_wmask,
  input  [63:0] io_rw_req_bits_wdata,
  input         io_rw_resp_ready,
  output        io_rw_resp_valid,
  output [63:0] io_rw_resp_bits_rdata,
  output        io_difftestCtrl_enable,
  output        io_meip,
  input         io_dma_aw_ready,
  output        io_dma_aw_valid,
  output [31:0] io_dma_aw_bits_addr,
  output [7:0]  io_dma_aw_bits_len,
  output [2:0]  io_dma_aw_bits_size,
  input         io_dma_w_ready,
  output        io_dma_w_valid,
  output [63:0] io_dma_w_bits_data,
  output [7:0]  io_dma_w_bits_strb,
  output        io_dma_b_ready,
  input         io_dma_b_valid,
  input         io_dma_ar_ready,
  output        io_dma_ar_valid,
  output [31:0] io_dma_ar_bits_addr,
  output        io_dma_r_ready,
  input         io_dma_r_valid,
  input  [63:0] io_dma_r_bits_data,
  input         _T_13
);
  wire  xbar_clock; // @[SimMMIO.scala 45:20]
  wire  xbar_reset; // @[SimMMIO.scala 45:20]
  wire  xbar_io_in_req_ready; // @[SimMMIO.scala 45:20]
  wire  xbar_io_in_req_valid; // @[SimMMIO.scala 45:20]
  wire [31:0] xbar_io_in_req_bits_addr; // @[SimMMIO.scala 45:20]
  wire [2:0] xbar_io_in_req_bits_size; // @[SimMMIO.scala 45:20]
  wire [3:0] xbar_io_in_req_bits_cmd; // @[SimMMIO.scala 45:20]
  wire [7:0] xbar_io_in_req_bits_wmask; // @[SimMMIO.scala 45:20]
  wire [63:0] xbar_io_in_req_bits_wdata; // @[SimMMIO.scala 45:20]
  wire  xbar_io_in_resp_ready; // @[SimMMIO.scala 45:20]
  wire  xbar_io_in_resp_valid; // @[SimMMIO.scala 45:20]
  wire [3:0] xbar_io_in_resp_bits_cmd; // @[SimMMIO.scala 45:20]
  wire [63:0] xbar_io_in_resp_bits_rdata; // @[SimMMIO.scala 45:20]
  wire  xbar_io_out_0_req_ready; // @[SimMMIO.scala 45:20]
  wire  xbar_io_out_0_req_valid; // @[SimMMIO.scala 45:20]
  wire [31:0] xbar_io_out_0_req_bits_addr; // @[SimMMIO.scala 45:20]
  wire [2:0] xbar_io_out_0_req_bits_size; // @[SimMMIO.scala 45:20]
  wire [3:0] xbar_io_out_0_req_bits_cmd; // @[SimMMIO.scala 45:20]
  wire [7:0] xbar_io_out_0_req_bits_wmask; // @[SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_0_req_bits_wdata; // @[SimMMIO.scala 45:20]
  wire  xbar_io_out_0_resp_ready; // @[SimMMIO.scala 45:20]
  wire  xbar_io_out_0_resp_valid; // @[SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_0_resp_bits_rdata; // @[SimMMIO.scala 45:20]
  wire  xbar_io_out_1_req_ready; // @[SimMMIO.scala 45:20]
  wire  xbar_io_out_1_req_valid; // @[SimMMIO.scala 45:20]
  wire [31:0] xbar_io_out_1_req_bits_addr; // @[SimMMIO.scala 45:20]
  wire [2:0] xbar_io_out_1_req_bits_size; // @[SimMMIO.scala 45:20]
  wire [3:0] xbar_io_out_1_req_bits_cmd; // @[SimMMIO.scala 45:20]
  wire [7:0] xbar_io_out_1_req_bits_wmask; // @[SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_1_req_bits_wdata; // @[SimMMIO.scala 45:20]
  wire  xbar_io_out_1_resp_ready; // @[SimMMIO.scala 45:20]
  wire  xbar_io_out_1_resp_valid; // @[SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_1_resp_bits_rdata; // @[SimMMIO.scala 45:20]
  wire  xbar_io_out_2_req_ready; // @[SimMMIO.scala 45:20]
  wire  xbar_io_out_2_req_valid; // @[SimMMIO.scala 45:20]
  wire [31:0] xbar_io_out_2_req_bits_addr; // @[SimMMIO.scala 45:20]
  wire [2:0] xbar_io_out_2_req_bits_size; // @[SimMMIO.scala 45:20]
  wire [3:0] xbar_io_out_2_req_bits_cmd; // @[SimMMIO.scala 45:20]
  wire [7:0] xbar_io_out_2_req_bits_wmask; // @[SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_2_req_bits_wdata; // @[SimMMIO.scala 45:20]
  wire  xbar_io_out_2_resp_ready; // @[SimMMIO.scala 45:20]
  wire  xbar_io_out_2_resp_valid; // @[SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_2_resp_bits_rdata; // @[SimMMIO.scala 45:20]
  wire  xbar_io_out_3_req_ready; // @[SimMMIO.scala 45:20]
  wire  xbar_io_out_3_req_valid; // @[SimMMIO.scala 45:20]
  wire [31:0] xbar_io_out_3_req_bits_addr; // @[SimMMIO.scala 45:20]
  wire [2:0] xbar_io_out_3_req_bits_size; // @[SimMMIO.scala 45:20]
  wire [3:0] xbar_io_out_3_req_bits_cmd; // @[SimMMIO.scala 45:20]
  wire [7:0] xbar_io_out_3_req_bits_wmask; // @[SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_3_req_bits_wdata; // @[SimMMIO.scala 45:20]
  wire  xbar_io_out_3_resp_ready; // @[SimMMIO.scala 45:20]
  wire  xbar_io_out_3_resp_valid; // @[SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_3_resp_bits_rdata; // @[SimMMIO.scala 45:20]
  wire  xbar_io_out_4_req_ready; // @[SimMMIO.scala 45:20]
  wire  xbar_io_out_4_req_valid; // @[SimMMIO.scala 45:20]
  wire [31:0] xbar_io_out_4_req_bits_addr; // @[SimMMIO.scala 45:20]
  wire [2:0] xbar_io_out_4_req_bits_size; // @[SimMMIO.scala 45:20]
  wire [3:0] xbar_io_out_4_req_bits_cmd; // @[SimMMIO.scala 45:20]
  wire [7:0] xbar_io_out_4_req_bits_wmask; // @[SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_4_req_bits_wdata; // @[SimMMIO.scala 45:20]
  wire  xbar_io_out_4_resp_ready; // @[SimMMIO.scala 45:20]
  wire  xbar_io_out_4_resp_valid; // @[SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_4_resp_bits_rdata; // @[SimMMIO.scala 45:20]
  wire  xbar_io_out_5_req_ready; // @[SimMMIO.scala 45:20]
  wire  xbar_io_out_5_req_valid; // @[SimMMIO.scala 45:20]
  wire [31:0] xbar_io_out_5_req_bits_addr; // @[SimMMIO.scala 45:20]
  wire [2:0] xbar_io_out_5_req_bits_size; // @[SimMMIO.scala 45:20]
  wire [3:0] xbar_io_out_5_req_bits_cmd; // @[SimMMIO.scala 45:20]
  wire [7:0] xbar_io_out_5_req_bits_wmask; // @[SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_5_req_bits_wdata; // @[SimMMIO.scala 45:20]
  wire  xbar_io_out_5_resp_ready; // @[SimMMIO.scala 45:20]
  wire  xbar_io_out_5_resp_valid; // @[SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_5_resp_bits_rdata; // @[SimMMIO.scala 45:20]
  wire  xbar_io_out_6_req_ready; // @[SimMMIO.scala 45:20]
  wire  xbar_io_out_6_req_valid; // @[SimMMIO.scala 45:20]
  wire [31:0] xbar_io_out_6_req_bits_addr; // @[SimMMIO.scala 45:20]
  wire [2:0] xbar_io_out_6_req_bits_size; // @[SimMMIO.scala 45:20]
  wire [3:0] xbar_io_out_6_req_bits_cmd; // @[SimMMIO.scala 45:20]
  wire [7:0] xbar_io_out_6_req_bits_wmask; // @[SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_6_req_bits_wdata; // @[SimMMIO.scala 45:20]
  wire  xbar_io_out_6_resp_ready; // @[SimMMIO.scala 45:20]
  wire  xbar_io_out_6_resp_valid; // @[SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_6_resp_bits_rdata; // @[SimMMIO.scala 45:20]
  wire  xbar_io_out_7_req_ready; // @[SimMMIO.scala 45:20]
  wire  xbar_io_out_7_req_valid; // @[SimMMIO.scala 45:20]
  wire [31:0] xbar_io_out_7_req_bits_addr; // @[SimMMIO.scala 45:20]
  wire [2:0] xbar_io_out_7_req_bits_size; // @[SimMMIO.scala 45:20]
  wire [3:0] xbar_io_out_7_req_bits_cmd; // @[SimMMIO.scala 45:20]
  wire [7:0] xbar_io_out_7_req_bits_wmask; // @[SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_7_req_bits_wdata; // @[SimMMIO.scala 45:20]
  wire  xbar_io_out_7_resp_ready; // @[SimMMIO.scala 45:20]
  wire  xbar_io_out_7_resp_valid; // @[SimMMIO.scala 45:20]
  wire [63:0] xbar_io_out_7_resp_bits_rdata; // @[SimMMIO.scala 45:20]
  wire  xbar_DISPLAY_ENABLE; // @[SimMMIO.scala 45:20]
  wire  uart_clock; // @[SimMMIO.scala 48:20]
  wire  uart_reset; // @[SimMMIO.scala 48:20]
  wire  uart_io_in_aw_ready; // @[SimMMIO.scala 48:20]
  wire  uart_io_in_aw_valid; // @[SimMMIO.scala 48:20]
  wire [31:0] uart_io_in_aw_bits_addr; // @[SimMMIO.scala 48:20]
  wire  uart_io_in_w_ready; // @[SimMMIO.scala 48:20]
  wire  uart_io_in_w_valid; // @[SimMMIO.scala 48:20]
  wire [63:0] uart_io_in_w_bits_data; // @[SimMMIO.scala 48:20]
  wire [7:0] uart_io_in_w_bits_strb; // @[SimMMIO.scala 48:20]
  wire  uart_io_in_b_ready; // @[SimMMIO.scala 48:20]
  wire  uart_io_in_b_valid; // @[SimMMIO.scala 48:20]
  wire  uart_io_in_ar_ready; // @[SimMMIO.scala 48:20]
  wire  uart_io_in_ar_valid; // @[SimMMIO.scala 48:20]
  wire [31:0] uart_io_in_ar_bits_addr; // @[SimMMIO.scala 48:20]
  wire  uart_io_in_r_ready; // @[SimMMIO.scala 48:20]
  wire  uart_io_in_r_valid; // @[SimMMIO.scala 48:20]
  wire [63:0] uart_io_in_r_bits_data; // @[SimMMIO.scala 48:20]
  wire  vga_clock; // @[SimMMIO.scala 49:19]
  wire  vga_reset; // @[SimMMIO.scala 49:19]
  wire  vga_io_in_fb_aw_ready; // @[SimMMIO.scala 49:19]
  wire  vga_io_in_fb_aw_valid; // @[SimMMIO.scala 49:19]
  wire [31:0] vga_io_in_fb_aw_bits_addr; // @[SimMMIO.scala 49:19]
  wire  vga_io_in_fb_w_ready; // @[SimMMIO.scala 49:19]
  wire  vga_io_in_fb_w_valid; // @[SimMMIO.scala 49:19]
  wire [63:0] vga_io_in_fb_w_bits_data; // @[SimMMIO.scala 49:19]
  wire [7:0] vga_io_in_fb_w_bits_strb; // @[SimMMIO.scala 49:19]
  wire  vga_io_in_fb_b_ready; // @[SimMMIO.scala 49:19]
  wire  vga_io_in_fb_b_valid; // @[SimMMIO.scala 49:19]
  wire  vga_io_in_fb_ar_ready; // @[SimMMIO.scala 49:19]
  wire  vga_io_in_fb_ar_valid; // @[SimMMIO.scala 49:19]
  wire  vga_io_in_fb_r_ready; // @[SimMMIO.scala 49:19]
  wire  vga_io_in_fb_r_valid; // @[SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_aw_ready; // @[SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_aw_valid; // @[SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_w_ready; // @[SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_w_valid; // @[SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_b_ready; // @[SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_b_valid; // @[SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_ar_ready; // @[SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_ar_valid; // @[SimMMIO.scala 49:19]
  wire [31:0] vga_io_in_ctrl_ar_bits_addr; // @[SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_r_ready; // @[SimMMIO.scala 49:19]
  wire  vga_io_in_ctrl_r_valid; // @[SimMMIO.scala 49:19]
  wire [63:0] vga_io_in_ctrl_r_bits_data; // @[SimMMIO.scala 49:19]
  wire  vga_io_vga_valid; // @[SimMMIO.scala 49:19]
  wire  flash_clock; // @[SimMMIO.scala 50:21]
  wire  flash_reset; // @[SimMMIO.scala 50:21]
  wire  flash_io_in_aw_ready; // @[SimMMIO.scala 50:21]
  wire  flash_io_in_aw_valid; // @[SimMMIO.scala 50:21]
  wire  flash_io_in_w_ready; // @[SimMMIO.scala 50:21]
  wire  flash_io_in_w_valid; // @[SimMMIO.scala 50:21]
  wire  flash_io_in_b_ready; // @[SimMMIO.scala 50:21]
  wire  flash_io_in_b_valid; // @[SimMMIO.scala 50:21]
  wire  flash_io_in_ar_ready; // @[SimMMIO.scala 50:21]
  wire  flash_io_in_ar_valid; // @[SimMMIO.scala 50:21]
  wire [31:0] flash_io_in_ar_bits_addr; // @[SimMMIO.scala 50:21]
  wire  flash_io_in_r_ready; // @[SimMMIO.scala 50:21]
  wire  flash_io_in_r_valid; // @[SimMMIO.scala 50:21]
  wire [63:0] flash_io_in_r_bits_data; // @[SimMMIO.scala 50:21]
  wire  sd_clock; // @[SimMMIO.scala 51:18]
  wire  sd_reset; // @[SimMMIO.scala 51:18]
  wire  sd_io_in_aw_ready; // @[SimMMIO.scala 51:18]
  wire  sd_io_in_aw_valid; // @[SimMMIO.scala 51:18]
  wire [31:0] sd_io_in_aw_bits_addr; // @[SimMMIO.scala 51:18]
  wire  sd_io_in_w_ready; // @[SimMMIO.scala 51:18]
  wire  sd_io_in_w_valid; // @[SimMMIO.scala 51:18]
  wire [63:0] sd_io_in_w_bits_data; // @[SimMMIO.scala 51:18]
  wire [7:0] sd_io_in_w_bits_strb; // @[SimMMIO.scala 51:18]
  wire  sd_io_in_b_ready; // @[SimMMIO.scala 51:18]
  wire  sd_io_in_b_valid; // @[SimMMIO.scala 51:18]
  wire  sd_io_in_ar_ready; // @[SimMMIO.scala 51:18]
  wire  sd_io_in_ar_valid; // @[SimMMIO.scala 51:18]
  wire [31:0] sd_io_in_ar_bits_addr; // @[SimMMIO.scala 51:18]
  wire  sd_io_in_r_ready; // @[SimMMIO.scala 51:18]
  wire  sd_io_in_r_valid; // @[SimMMIO.scala 51:18]
  wire [63:0] sd_io_in_r_bits_data; // @[SimMMIO.scala 51:18]
  wire  difftestCtrl_clock; // @[SimMMIO.scala 52:28]
  wire  difftestCtrl_reset; // @[SimMMIO.scala 52:28]
  wire  difftestCtrl_io_in_aw_ready; // @[SimMMIO.scala 52:28]
  wire  difftestCtrl_io_in_aw_valid; // @[SimMMIO.scala 52:28]
  wire [31:0] difftestCtrl_io_in_aw_bits_addr; // @[SimMMIO.scala 52:28]
  wire  difftestCtrl_io_in_w_ready; // @[SimMMIO.scala 52:28]
  wire  difftestCtrl_io_in_w_valid; // @[SimMMIO.scala 52:28]
  wire [63:0] difftestCtrl_io_in_w_bits_data; // @[SimMMIO.scala 52:28]
  wire [7:0] difftestCtrl_io_in_w_bits_strb; // @[SimMMIO.scala 52:28]
  wire  difftestCtrl_io_in_b_ready; // @[SimMMIO.scala 52:28]
  wire  difftestCtrl_io_in_b_valid; // @[SimMMIO.scala 52:28]
  wire  difftestCtrl_io_in_ar_ready; // @[SimMMIO.scala 52:28]
  wire  difftestCtrl_io_in_ar_valid; // @[SimMMIO.scala 52:28]
  wire  difftestCtrl_io_in_r_ready; // @[SimMMIO.scala 52:28]
  wire  difftestCtrl_io_in_r_valid; // @[SimMMIO.scala 52:28]
  wire [63:0] difftestCtrl_io_in_r_bits_data; // @[SimMMIO.scala 52:28]
  wire  difftestCtrl_io_extra_enable; // @[SimMMIO.scala 52:28]
  wire  meipGen_clock; // @[SimMMIO.scala 53:23]
  wire  meipGen_reset; // @[SimMMIO.scala 53:23]
  wire  meipGen_io_in_aw_ready; // @[SimMMIO.scala 53:23]
  wire  meipGen_io_in_aw_valid; // @[SimMMIO.scala 53:23]
  wire [31:0] meipGen_io_in_aw_bits_addr; // @[SimMMIO.scala 53:23]
  wire  meipGen_io_in_w_ready; // @[SimMMIO.scala 53:23]
  wire  meipGen_io_in_w_valid; // @[SimMMIO.scala 53:23]
  wire [63:0] meipGen_io_in_w_bits_data; // @[SimMMIO.scala 53:23]
  wire [7:0] meipGen_io_in_w_bits_strb; // @[SimMMIO.scala 53:23]
  wire  meipGen_io_in_b_ready; // @[SimMMIO.scala 53:23]
  wire  meipGen_io_in_b_valid; // @[SimMMIO.scala 53:23]
  wire  meipGen_io_in_ar_ready; // @[SimMMIO.scala 53:23]
  wire  meipGen_io_in_ar_valid; // @[SimMMIO.scala 53:23]
  wire  meipGen_io_in_r_ready; // @[SimMMIO.scala 53:23]
  wire  meipGen_io_in_r_valid; // @[SimMMIO.scala 53:23]
  wire [63:0] meipGen_io_in_r_bits_data; // @[SimMMIO.scala 53:23]
  wire  meipGen_io_extra_enable; // @[SimMMIO.scala 53:23]
  wire  dma_clock; // @[SimMMIO.scala 54:19]
  wire  dma_reset; // @[SimMMIO.scala 54:19]
  wire  dma_io_in_aw_ready; // @[SimMMIO.scala 54:19]
  wire  dma_io_in_aw_valid; // @[SimMMIO.scala 54:19]
  wire [31:0] dma_io_in_aw_bits_addr; // @[SimMMIO.scala 54:19]
  wire  dma_io_in_w_ready; // @[SimMMIO.scala 54:19]
  wire  dma_io_in_w_valid; // @[SimMMIO.scala 54:19]
  wire [63:0] dma_io_in_w_bits_data; // @[SimMMIO.scala 54:19]
  wire [7:0] dma_io_in_w_bits_strb; // @[SimMMIO.scala 54:19]
  wire  dma_io_in_b_ready; // @[SimMMIO.scala 54:19]
  wire  dma_io_in_b_valid; // @[SimMMIO.scala 54:19]
  wire  dma_io_in_ar_ready; // @[SimMMIO.scala 54:19]
  wire  dma_io_in_ar_valid; // @[SimMMIO.scala 54:19]
  wire [31:0] dma_io_in_ar_bits_addr; // @[SimMMIO.scala 54:19]
  wire  dma_io_in_r_ready; // @[SimMMIO.scala 54:19]
  wire  dma_io_in_r_valid; // @[SimMMIO.scala 54:19]
  wire [63:0] dma_io_in_r_bits_data; // @[SimMMIO.scala 54:19]
  wire  dma_io_extra_dma_aw_ready; // @[SimMMIO.scala 54:19]
  wire  dma_io_extra_dma_aw_valid; // @[SimMMIO.scala 54:19]
  wire [31:0] dma_io_extra_dma_aw_bits_addr; // @[SimMMIO.scala 54:19]
  wire [7:0] dma_io_extra_dma_aw_bits_len; // @[SimMMIO.scala 54:19]
  wire [2:0] dma_io_extra_dma_aw_bits_size; // @[SimMMIO.scala 54:19]
  wire  dma_io_extra_dma_w_ready; // @[SimMMIO.scala 54:19]
  wire  dma_io_extra_dma_w_valid; // @[SimMMIO.scala 54:19]
  wire [63:0] dma_io_extra_dma_w_bits_data; // @[SimMMIO.scala 54:19]
  wire [7:0] dma_io_extra_dma_w_bits_strb; // @[SimMMIO.scala 54:19]
  wire  dma_io_extra_dma_w_bits_last; // @[SimMMIO.scala 54:19]
  wire  dma_io_extra_dma_b_ready; // @[SimMMIO.scala 54:19]
  wire  dma_io_extra_dma_b_valid; // @[SimMMIO.scala 54:19]
  wire  dma_io_extra_dma_ar_ready; // @[SimMMIO.scala 54:19]
  wire  dma_io_extra_dma_ar_valid; // @[SimMMIO.scala 54:19]
  wire [31:0] dma_io_extra_dma_ar_bits_addr; // @[SimMMIO.scala 54:19]
  wire [7:0] dma_io_extra_dma_ar_bits_len; // @[SimMMIO.scala 54:19]
  wire [2:0] dma_io_extra_dma_ar_bits_size; // @[SimMMIO.scala 54:19]
  wire  dma_io_extra_dma_r_ready; // @[SimMMIO.scala 54:19]
  wire  dma_io_extra_dma_r_valid; // @[SimMMIO.scala 54:19]
  wire [63:0] dma_io_extra_dma_r_bits_data; // @[SimMMIO.scala 54:19]
  wire  SimpleBus2AXI4Converter_clock; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_reset; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_in_req_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_in_req_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_io_in_req_bits_addr; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_io_in_req_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_io_in_req_bits_wmask; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_io_in_req_bits_wdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_in_resp_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_in_resp_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_io_in_resp_bits_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_aw_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_aw_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_io_out_aw_bits_addr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_w_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_w_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_io_out_w_bits_data; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_io_out_w_bits_strb; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_b_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_b_valid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_ar_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_ar_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_io_out_ar_bits_addr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_r_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_r_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_io_out_r_bits_data; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_clock; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_reset; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_in_req_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_in_req_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_1_io_in_req_bits_addr; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_1_io_in_req_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_1_io_in_req_bits_wmask; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_1_io_in_req_bits_wdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_in_resp_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_in_resp_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_1_io_in_resp_bits_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_aw_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_aw_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_1_io_out_aw_bits_addr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_w_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_w_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_1_io_out_w_bits_data; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_1_io_out_w_bits_strb; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_b_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_b_valid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_ar_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_ar_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_1_io_out_ar_bits_addr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_r_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_r_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_1_io_out_r_bits_data; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_clock; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_reset; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_in_req_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_in_req_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_2_io_in_req_bits_addr; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_2_io_in_req_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_2_io_in_req_bits_wmask; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_2_io_in_req_bits_wdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_in_resp_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_in_resp_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_2_io_in_resp_bits_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_aw_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_aw_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_2_io_out_aw_bits_addr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_w_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_w_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_2_io_out_w_bits_data; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_2_io_out_w_bits_strb; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_b_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_b_valid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_ar_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_ar_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_2_io_out_ar_bits_addr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_r_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_r_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_2_io_out_r_bits_data; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_clock; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_reset; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_in_req_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_in_req_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_3_io_in_req_bits_addr; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_3_io_in_req_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_3_io_in_req_bits_wmask; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_3_io_in_req_bits_wdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_in_resp_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_in_resp_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_3_io_in_resp_bits_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_aw_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_aw_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_3_io_out_aw_bits_addr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_w_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_w_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_3_io_out_w_bits_data; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_3_io_out_w_bits_strb; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_b_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_b_valid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_ar_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_ar_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_3_io_out_ar_bits_addr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_r_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_r_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_3_io_out_r_bits_data; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_4_clock; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_4_reset; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_4_io_in_req_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_4_io_in_req_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_4_io_in_req_bits_addr; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_4_io_in_req_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_4_io_in_req_bits_wmask; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_4_io_in_req_bits_wdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_4_io_in_resp_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_4_io_in_resp_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_4_io_in_resp_bits_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_4_io_out_aw_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_4_io_out_aw_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_4_io_out_aw_bits_addr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_4_io_out_w_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_4_io_out_w_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_4_io_out_w_bits_data; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_4_io_out_w_bits_strb; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_4_io_out_b_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_4_io_out_b_valid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_4_io_out_ar_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_4_io_out_ar_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_4_io_out_ar_bits_addr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_4_io_out_r_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_4_io_out_r_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_4_io_out_r_bits_data; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_5_clock; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_5_reset; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_5_io_in_req_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_5_io_in_req_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_5_io_in_req_bits_addr; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_5_io_in_req_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_5_io_in_req_bits_wmask; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_5_io_in_req_bits_wdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_5_io_in_resp_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_5_io_in_resp_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_5_io_in_resp_bits_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_5_io_out_aw_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_5_io_out_aw_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_5_io_out_aw_bits_addr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_5_io_out_w_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_5_io_out_w_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_5_io_out_w_bits_data; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_5_io_out_w_bits_strb; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_5_io_out_b_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_5_io_out_b_valid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_5_io_out_ar_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_5_io_out_ar_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_5_io_out_ar_bits_addr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_5_io_out_r_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_5_io_out_r_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_5_io_out_r_bits_data; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_6_clock; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_6_reset; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_6_io_in_req_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_6_io_in_req_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_6_io_in_req_bits_addr; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_6_io_in_req_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_6_io_in_req_bits_wmask; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_6_io_in_req_bits_wdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_6_io_in_resp_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_6_io_in_resp_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_6_io_in_resp_bits_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_6_io_out_aw_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_6_io_out_aw_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_6_io_out_aw_bits_addr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_6_io_out_w_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_6_io_out_w_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_6_io_out_w_bits_data; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_6_io_out_w_bits_strb; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_6_io_out_b_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_6_io_out_b_valid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_6_io_out_ar_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_6_io_out_ar_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_6_io_out_ar_bits_addr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_6_io_out_r_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_6_io_out_r_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_6_io_out_r_bits_data; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_7_clock; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_7_reset; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_7_io_in_req_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_7_io_in_req_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_7_io_in_req_bits_addr; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_7_io_in_req_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_7_io_in_req_bits_wmask; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_7_io_in_req_bits_wdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_7_io_in_resp_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_7_io_in_resp_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_7_io_in_resp_bits_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_7_io_out_aw_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_7_io_out_aw_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_7_io_out_aw_bits_addr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_7_io_out_w_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_7_io_out_w_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_7_io_out_w_bits_data; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_7_io_out_w_bits_strb; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_7_io_out_b_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_7_io_out_b_valid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_7_io_out_ar_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_7_io_out_ar_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_7_io_out_ar_bits_addr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_7_io_out_r_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_7_io_out_r_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_7_io_out_r_bits_data; // @[ToAXI4.scala 204:24]
  SimpleBusCrossbar1toN_1 xbar ( // @[SimMMIO.scala 45:20]
    .clock(xbar_clock),
    .reset(xbar_reset),
    .io_in_req_ready(xbar_io_in_req_ready),
    .io_in_req_valid(xbar_io_in_req_valid),
    .io_in_req_bits_addr(xbar_io_in_req_bits_addr),
    .io_in_req_bits_size(xbar_io_in_req_bits_size),
    .io_in_req_bits_cmd(xbar_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(xbar_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(xbar_io_in_req_bits_wdata),
    .io_in_resp_ready(xbar_io_in_resp_ready),
    .io_in_resp_valid(xbar_io_in_resp_valid),
    .io_in_resp_bits_cmd(xbar_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(xbar_io_in_resp_bits_rdata),
    .io_out_0_req_ready(xbar_io_out_0_req_ready),
    .io_out_0_req_valid(xbar_io_out_0_req_valid),
    .io_out_0_req_bits_addr(xbar_io_out_0_req_bits_addr),
    .io_out_0_req_bits_size(xbar_io_out_0_req_bits_size),
    .io_out_0_req_bits_cmd(xbar_io_out_0_req_bits_cmd),
    .io_out_0_req_bits_wmask(xbar_io_out_0_req_bits_wmask),
    .io_out_0_req_bits_wdata(xbar_io_out_0_req_bits_wdata),
    .io_out_0_resp_ready(xbar_io_out_0_resp_ready),
    .io_out_0_resp_valid(xbar_io_out_0_resp_valid),
    .io_out_0_resp_bits_rdata(xbar_io_out_0_resp_bits_rdata),
    .io_out_1_req_ready(xbar_io_out_1_req_ready),
    .io_out_1_req_valid(xbar_io_out_1_req_valid),
    .io_out_1_req_bits_addr(xbar_io_out_1_req_bits_addr),
    .io_out_1_req_bits_size(xbar_io_out_1_req_bits_size),
    .io_out_1_req_bits_cmd(xbar_io_out_1_req_bits_cmd),
    .io_out_1_req_bits_wmask(xbar_io_out_1_req_bits_wmask),
    .io_out_1_req_bits_wdata(xbar_io_out_1_req_bits_wdata),
    .io_out_1_resp_ready(xbar_io_out_1_resp_ready),
    .io_out_1_resp_valid(xbar_io_out_1_resp_valid),
    .io_out_1_resp_bits_rdata(xbar_io_out_1_resp_bits_rdata),
    .io_out_2_req_ready(xbar_io_out_2_req_ready),
    .io_out_2_req_valid(xbar_io_out_2_req_valid),
    .io_out_2_req_bits_addr(xbar_io_out_2_req_bits_addr),
    .io_out_2_req_bits_size(xbar_io_out_2_req_bits_size),
    .io_out_2_req_bits_cmd(xbar_io_out_2_req_bits_cmd),
    .io_out_2_req_bits_wmask(xbar_io_out_2_req_bits_wmask),
    .io_out_2_req_bits_wdata(xbar_io_out_2_req_bits_wdata),
    .io_out_2_resp_ready(xbar_io_out_2_resp_ready),
    .io_out_2_resp_valid(xbar_io_out_2_resp_valid),
    .io_out_2_resp_bits_rdata(xbar_io_out_2_resp_bits_rdata),
    .io_out_3_req_ready(xbar_io_out_3_req_ready),
    .io_out_3_req_valid(xbar_io_out_3_req_valid),
    .io_out_3_req_bits_addr(xbar_io_out_3_req_bits_addr),
    .io_out_3_req_bits_size(xbar_io_out_3_req_bits_size),
    .io_out_3_req_bits_cmd(xbar_io_out_3_req_bits_cmd),
    .io_out_3_req_bits_wmask(xbar_io_out_3_req_bits_wmask),
    .io_out_3_req_bits_wdata(xbar_io_out_3_req_bits_wdata),
    .io_out_3_resp_ready(xbar_io_out_3_resp_ready),
    .io_out_3_resp_valid(xbar_io_out_3_resp_valid),
    .io_out_3_resp_bits_rdata(xbar_io_out_3_resp_bits_rdata),
    .io_out_4_req_ready(xbar_io_out_4_req_ready),
    .io_out_4_req_valid(xbar_io_out_4_req_valid),
    .io_out_4_req_bits_addr(xbar_io_out_4_req_bits_addr),
    .io_out_4_req_bits_size(xbar_io_out_4_req_bits_size),
    .io_out_4_req_bits_cmd(xbar_io_out_4_req_bits_cmd),
    .io_out_4_req_bits_wmask(xbar_io_out_4_req_bits_wmask),
    .io_out_4_req_bits_wdata(xbar_io_out_4_req_bits_wdata),
    .io_out_4_resp_ready(xbar_io_out_4_resp_ready),
    .io_out_4_resp_valid(xbar_io_out_4_resp_valid),
    .io_out_4_resp_bits_rdata(xbar_io_out_4_resp_bits_rdata),
    .io_out_5_req_ready(xbar_io_out_5_req_ready),
    .io_out_5_req_valid(xbar_io_out_5_req_valid),
    .io_out_5_req_bits_addr(xbar_io_out_5_req_bits_addr),
    .io_out_5_req_bits_size(xbar_io_out_5_req_bits_size),
    .io_out_5_req_bits_cmd(xbar_io_out_5_req_bits_cmd),
    .io_out_5_req_bits_wmask(xbar_io_out_5_req_bits_wmask),
    .io_out_5_req_bits_wdata(xbar_io_out_5_req_bits_wdata),
    .io_out_5_resp_ready(xbar_io_out_5_resp_ready),
    .io_out_5_resp_valid(xbar_io_out_5_resp_valid),
    .io_out_5_resp_bits_rdata(xbar_io_out_5_resp_bits_rdata),
    .io_out_6_req_ready(xbar_io_out_6_req_ready),
    .io_out_6_req_valid(xbar_io_out_6_req_valid),
    .io_out_6_req_bits_addr(xbar_io_out_6_req_bits_addr),
    .io_out_6_req_bits_size(xbar_io_out_6_req_bits_size),
    .io_out_6_req_bits_cmd(xbar_io_out_6_req_bits_cmd),
    .io_out_6_req_bits_wmask(xbar_io_out_6_req_bits_wmask),
    .io_out_6_req_bits_wdata(xbar_io_out_6_req_bits_wdata),
    .io_out_6_resp_ready(xbar_io_out_6_resp_ready),
    .io_out_6_resp_valid(xbar_io_out_6_resp_valid),
    .io_out_6_resp_bits_rdata(xbar_io_out_6_resp_bits_rdata),
    .io_out_7_req_ready(xbar_io_out_7_req_ready),
    .io_out_7_req_valid(xbar_io_out_7_req_valid),
    .io_out_7_req_bits_addr(xbar_io_out_7_req_bits_addr),
    .io_out_7_req_bits_size(xbar_io_out_7_req_bits_size),
    .io_out_7_req_bits_cmd(xbar_io_out_7_req_bits_cmd),
    .io_out_7_req_bits_wmask(xbar_io_out_7_req_bits_wmask),
    .io_out_7_req_bits_wdata(xbar_io_out_7_req_bits_wdata),
    .io_out_7_resp_ready(xbar_io_out_7_resp_ready),
    .io_out_7_resp_valid(xbar_io_out_7_resp_valid),
    .io_out_7_resp_bits_rdata(xbar_io_out_7_resp_bits_rdata),
    .DISPLAY_ENABLE(xbar_DISPLAY_ENABLE)
  );
  AXI4UART uart ( // @[SimMMIO.scala 48:20]
    .clock(uart_clock),
    .reset(uart_reset),
    .io_in_aw_ready(uart_io_in_aw_ready),
    .io_in_aw_valid(uart_io_in_aw_valid),
    .io_in_aw_bits_addr(uart_io_in_aw_bits_addr),
    .io_in_w_ready(uart_io_in_w_ready),
    .io_in_w_valid(uart_io_in_w_valid),
    .io_in_w_bits_data(uart_io_in_w_bits_data),
    .io_in_w_bits_strb(uart_io_in_w_bits_strb),
    .io_in_b_ready(uart_io_in_b_ready),
    .io_in_b_valid(uart_io_in_b_valid),
    .io_in_ar_ready(uart_io_in_ar_ready),
    .io_in_ar_valid(uart_io_in_ar_valid),
    .io_in_ar_bits_addr(uart_io_in_ar_bits_addr),
    .io_in_r_ready(uart_io_in_r_ready),
    .io_in_r_valid(uart_io_in_r_valid),
    .io_in_r_bits_data(uart_io_in_r_bits_data)
  );
  AXI4VGA vga ( // @[SimMMIO.scala 49:19]
    .clock(vga_clock),
    .reset(vga_reset),
    .io_in_fb_aw_ready(vga_io_in_fb_aw_ready),
    .io_in_fb_aw_valid(vga_io_in_fb_aw_valid),
    .io_in_fb_aw_bits_addr(vga_io_in_fb_aw_bits_addr),
    .io_in_fb_w_ready(vga_io_in_fb_w_ready),
    .io_in_fb_w_valid(vga_io_in_fb_w_valid),
    .io_in_fb_w_bits_data(vga_io_in_fb_w_bits_data),
    .io_in_fb_w_bits_strb(vga_io_in_fb_w_bits_strb),
    .io_in_fb_b_ready(vga_io_in_fb_b_ready),
    .io_in_fb_b_valid(vga_io_in_fb_b_valid),
    .io_in_fb_ar_ready(vga_io_in_fb_ar_ready),
    .io_in_fb_ar_valid(vga_io_in_fb_ar_valid),
    .io_in_fb_r_ready(vga_io_in_fb_r_ready),
    .io_in_fb_r_valid(vga_io_in_fb_r_valid),
    .io_in_ctrl_aw_ready(vga_io_in_ctrl_aw_ready),
    .io_in_ctrl_aw_valid(vga_io_in_ctrl_aw_valid),
    .io_in_ctrl_w_ready(vga_io_in_ctrl_w_ready),
    .io_in_ctrl_w_valid(vga_io_in_ctrl_w_valid),
    .io_in_ctrl_b_ready(vga_io_in_ctrl_b_ready),
    .io_in_ctrl_b_valid(vga_io_in_ctrl_b_valid),
    .io_in_ctrl_ar_ready(vga_io_in_ctrl_ar_ready),
    .io_in_ctrl_ar_valid(vga_io_in_ctrl_ar_valid),
    .io_in_ctrl_ar_bits_addr(vga_io_in_ctrl_ar_bits_addr),
    .io_in_ctrl_r_ready(vga_io_in_ctrl_r_ready),
    .io_in_ctrl_r_valid(vga_io_in_ctrl_r_valid),
    .io_in_ctrl_r_bits_data(vga_io_in_ctrl_r_bits_data),
    .io_vga_valid(vga_io_vga_valid)
  );
  AXI4Flash flash ( // @[SimMMIO.scala 50:21]
    .clock(flash_clock),
    .reset(flash_reset),
    .io_in_aw_ready(flash_io_in_aw_ready),
    .io_in_aw_valid(flash_io_in_aw_valid),
    .io_in_w_ready(flash_io_in_w_ready),
    .io_in_w_valid(flash_io_in_w_valid),
    .io_in_b_ready(flash_io_in_b_ready),
    .io_in_b_valid(flash_io_in_b_valid),
    .io_in_ar_ready(flash_io_in_ar_ready),
    .io_in_ar_valid(flash_io_in_ar_valid),
    .io_in_ar_bits_addr(flash_io_in_ar_bits_addr),
    .io_in_r_ready(flash_io_in_r_ready),
    .io_in_r_valid(flash_io_in_r_valid),
    .io_in_r_bits_data(flash_io_in_r_bits_data)
  );
  AXI4DummySD sd ( // @[SimMMIO.scala 51:18]
    .clock(sd_clock),
    .reset(sd_reset),
    .io_in_aw_ready(sd_io_in_aw_ready),
    .io_in_aw_valid(sd_io_in_aw_valid),
    .io_in_aw_bits_addr(sd_io_in_aw_bits_addr),
    .io_in_w_ready(sd_io_in_w_ready),
    .io_in_w_valid(sd_io_in_w_valid),
    .io_in_w_bits_data(sd_io_in_w_bits_data),
    .io_in_w_bits_strb(sd_io_in_w_bits_strb),
    .io_in_b_ready(sd_io_in_b_ready),
    .io_in_b_valid(sd_io_in_b_valid),
    .io_in_ar_ready(sd_io_in_ar_ready),
    .io_in_ar_valid(sd_io_in_ar_valid),
    .io_in_ar_bits_addr(sd_io_in_ar_bits_addr),
    .io_in_r_ready(sd_io_in_r_ready),
    .io_in_r_valid(sd_io_in_r_valid),
    .io_in_r_bits_data(sd_io_in_r_bits_data)
  );
  AXI4DiffTestCtrl difftestCtrl ( // @[SimMMIO.scala 52:28]
    .clock(difftestCtrl_clock),
    .reset(difftestCtrl_reset),
    .io_in_aw_ready(difftestCtrl_io_in_aw_ready),
    .io_in_aw_valid(difftestCtrl_io_in_aw_valid),
    .io_in_aw_bits_addr(difftestCtrl_io_in_aw_bits_addr),
    .io_in_w_ready(difftestCtrl_io_in_w_ready),
    .io_in_w_valid(difftestCtrl_io_in_w_valid),
    .io_in_w_bits_data(difftestCtrl_io_in_w_bits_data),
    .io_in_w_bits_strb(difftestCtrl_io_in_w_bits_strb),
    .io_in_b_ready(difftestCtrl_io_in_b_ready),
    .io_in_b_valid(difftestCtrl_io_in_b_valid),
    .io_in_ar_ready(difftestCtrl_io_in_ar_ready),
    .io_in_ar_valid(difftestCtrl_io_in_ar_valid),
    .io_in_r_ready(difftestCtrl_io_in_r_ready),
    .io_in_r_valid(difftestCtrl_io_in_r_valid),
    .io_in_r_bits_data(difftestCtrl_io_in_r_bits_data),
    .io_extra_enable(difftestCtrl_io_extra_enable)
  );
  AXI4DiffTestCtrl meipGen ( // @[SimMMIO.scala 53:23]
    .clock(meipGen_clock),
    .reset(meipGen_reset),
    .io_in_aw_ready(meipGen_io_in_aw_ready),
    .io_in_aw_valid(meipGen_io_in_aw_valid),
    .io_in_aw_bits_addr(meipGen_io_in_aw_bits_addr),
    .io_in_w_ready(meipGen_io_in_w_ready),
    .io_in_w_valid(meipGen_io_in_w_valid),
    .io_in_w_bits_data(meipGen_io_in_w_bits_data),
    .io_in_w_bits_strb(meipGen_io_in_w_bits_strb),
    .io_in_b_ready(meipGen_io_in_b_ready),
    .io_in_b_valid(meipGen_io_in_b_valid),
    .io_in_ar_ready(meipGen_io_in_ar_ready),
    .io_in_ar_valid(meipGen_io_in_ar_valid),
    .io_in_r_ready(meipGen_io_in_r_ready),
    .io_in_r_valid(meipGen_io_in_r_valid),
    .io_in_r_bits_data(meipGen_io_in_r_bits_data),
    .io_extra_enable(meipGen_io_extra_enable)
  );
  AXI4DMA dma ( // @[SimMMIO.scala 54:19]
    .clock(dma_clock),
    .reset(dma_reset),
    .io_in_aw_ready(dma_io_in_aw_ready),
    .io_in_aw_valid(dma_io_in_aw_valid),
    .io_in_aw_bits_addr(dma_io_in_aw_bits_addr),
    .io_in_w_ready(dma_io_in_w_ready),
    .io_in_w_valid(dma_io_in_w_valid),
    .io_in_w_bits_data(dma_io_in_w_bits_data),
    .io_in_w_bits_strb(dma_io_in_w_bits_strb),
    .io_in_b_ready(dma_io_in_b_ready),
    .io_in_b_valid(dma_io_in_b_valid),
    .io_in_ar_ready(dma_io_in_ar_ready),
    .io_in_ar_valid(dma_io_in_ar_valid),
    .io_in_ar_bits_addr(dma_io_in_ar_bits_addr),
    .io_in_r_ready(dma_io_in_r_ready),
    .io_in_r_valid(dma_io_in_r_valid),
    .io_in_r_bits_data(dma_io_in_r_bits_data),
    .io_extra_dma_aw_ready(dma_io_extra_dma_aw_ready),
    .io_extra_dma_aw_valid(dma_io_extra_dma_aw_valid),
    .io_extra_dma_aw_bits_addr(dma_io_extra_dma_aw_bits_addr),
    .io_extra_dma_aw_bits_len(dma_io_extra_dma_aw_bits_len),
    .io_extra_dma_aw_bits_size(dma_io_extra_dma_aw_bits_size),
    .io_extra_dma_w_ready(dma_io_extra_dma_w_ready),
    .io_extra_dma_w_valid(dma_io_extra_dma_w_valid),
    .io_extra_dma_w_bits_data(dma_io_extra_dma_w_bits_data),
    .io_extra_dma_w_bits_strb(dma_io_extra_dma_w_bits_strb),
    .io_extra_dma_w_bits_last(dma_io_extra_dma_w_bits_last),
    .io_extra_dma_b_ready(dma_io_extra_dma_b_ready),
    .io_extra_dma_b_valid(dma_io_extra_dma_b_valid),
    .io_extra_dma_ar_ready(dma_io_extra_dma_ar_ready),
    .io_extra_dma_ar_valid(dma_io_extra_dma_ar_valid),
    .io_extra_dma_ar_bits_addr(dma_io_extra_dma_ar_bits_addr),
    .io_extra_dma_ar_bits_len(dma_io_extra_dma_ar_bits_len),
    .io_extra_dma_ar_bits_size(dma_io_extra_dma_ar_bits_size),
    .io_extra_dma_r_ready(dma_io_extra_dma_r_ready),
    .io_extra_dma_r_valid(dma_io_extra_dma_r_valid),
    .io_extra_dma_r_bits_data(dma_io_extra_dma_r_bits_data)
  );
  SimpleBus2AXI4Converter_1 SimpleBus2AXI4Converter ( // @[ToAXI4.scala 204:24]
    .clock(SimpleBus2AXI4Converter_clock),
    .reset(SimpleBus2AXI4Converter_reset),
    .io_in_req_ready(SimpleBus2AXI4Converter_io_in_req_ready),
    .io_in_req_valid(SimpleBus2AXI4Converter_io_in_req_valid),
    .io_in_req_bits_addr(SimpleBus2AXI4Converter_io_in_req_bits_addr),
    .io_in_req_bits_cmd(SimpleBus2AXI4Converter_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(SimpleBus2AXI4Converter_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(SimpleBus2AXI4Converter_io_in_req_bits_wdata),
    .io_in_resp_ready(SimpleBus2AXI4Converter_io_in_resp_ready),
    .io_in_resp_valid(SimpleBus2AXI4Converter_io_in_resp_valid),
    .io_in_resp_bits_rdata(SimpleBus2AXI4Converter_io_in_resp_bits_rdata),
    .io_out_aw_ready(SimpleBus2AXI4Converter_io_out_aw_ready),
    .io_out_aw_valid(SimpleBus2AXI4Converter_io_out_aw_valid),
    .io_out_aw_bits_addr(SimpleBus2AXI4Converter_io_out_aw_bits_addr),
    .io_out_w_ready(SimpleBus2AXI4Converter_io_out_w_ready),
    .io_out_w_valid(SimpleBus2AXI4Converter_io_out_w_valid),
    .io_out_w_bits_data(SimpleBus2AXI4Converter_io_out_w_bits_data),
    .io_out_w_bits_strb(SimpleBus2AXI4Converter_io_out_w_bits_strb),
    .io_out_b_ready(SimpleBus2AXI4Converter_io_out_b_ready),
    .io_out_b_valid(SimpleBus2AXI4Converter_io_out_b_valid),
    .io_out_ar_ready(SimpleBus2AXI4Converter_io_out_ar_ready),
    .io_out_ar_valid(SimpleBus2AXI4Converter_io_out_ar_valid),
    .io_out_ar_bits_addr(SimpleBus2AXI4Converter_io_out_ar_bits_addr),
    .io_out_r_ready(SimpleBus2AXI4Converter_io_out_r_ready),
    .io_out_r_valid(SimpleBus2AXI4Converter_io_out_r_valid),
    .io_out_r_bits_data(SimpleBus2AXI4Converter_io_out_r_bits_data)
  );
  SimpleBus2AXI4Converter_1 SimpleBus2AXI4Converter_1 ( // @[ToAXI4.scala 204:24]
    .clock(SimpleBus2AXI4Converter_1_clock),
    .reset(SimpleBus2AXI4Converter_1_reset),
    .io_in_req_ready(SimpleBus2AXI4Converter_1_io_in_req_ready),
    .io_in_req_valid(SimpleBus2AXI4Converter_1_io_in_req_valid),
    .io_in_req_bits_addr(SimpleBus2AXI4Converter_1_io_in_req_bits_addr),
    .io_in_req_bits_cmd(SimpleBus2AXI4Converter_1_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(SimpleBus2AXI4Converter_1_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(SimpleBus2AXI4Converter_1_io_in_req_bits_wdata),
    .io_in_resp_ready(SimpleBus2AXI4Converter_1_io_in_resp_ready),
    .io_in_resp_valid(SimpleBus2AXI4Converter_1_io_in_resp_valid),
    .io_in_resp_bits_rdata(SimpleBus2AXI4Converter_1_io_in_resp_bits_rdata),
    .io_out_aw_ready(SimpleBus2AXI4Converter_1_io_out_aw_ready),
    .io_out_aw_valid(SimpleBus2AXI4Converter_1_io_out_aw_valid),
    .io_out_aw_bits_addr(SimpleBus2AXI4Converter_1_io_out_aw_bits_addr),
    .io_out_w_ready(SimpleBus2AXI4Converter_1_io_out_w_ready),
    .io_out_w_valid(SimpleBus2AXI4Converter_1_io_out_w_valid),
    .io_out_w_bits_data(SimpleBus2AXI4Converter_1_io_out_w_bits_data),
    .io_out_w_bits_strb(SimpleBus2AXI4Converter_1_io_out_w_bits_strb),
    .io_out_b_ready(SimpleBus2AXI4Converter_1_io_out_b_ready),
    .io_out_b_valid(SimpleBus2AXI4Converter_1_io_out_b_valid),
    .io_out_ar_ready(SimpleBus2AXI4Converter_1_io_out_ar_ready),
    .io_out_ar_valid(SimpleBus2AXI4Converter_1_io_out_ar_valid),
    .io_out_ar_bits_addr(SimpleBus2AXI4Converter_1_io_out_ar_bits_addr),
    .io_out_r_ready(SimpleBus2AXI4Converter_1_io_out_r_ready),
    .io_out_r_valid(SimpleBus2AXI4Converter_1_io_out_r_valid),
    .io_out_r_bits_data(SimpleBus2AXI4Converter_1_io_out_r_bits_data)
  );
  SimpleBus2AXI4Converter_1 SimpleBus2AXI4Converter_2 ( // @[ToAXI4.scala 204:24]
    .clock(SimpleBus2AXI4Converter_2_clock),
    .reset(SimpleBus2AXI4Converter_2_reset),
    .io_in_req_ready(SimpleBus2AXI4Converter_2_io_in_req_ready),
    .io_in_req_valid(SimpleBus2AXI4Converter_2_io_in_req_valid),
    .io_in_req_bits_addr(SimpleBus2AXI4Converter_2_io_in_req_bits_addr),
    .io_in_req_bits_cmd(SimpleBus2AXI4Converter_2_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(SimpleBus2AXI4Converter_2_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(SimpleBus2AXI4Converter_2_io_in_req_bits_wdata),
    .io_in_resp_ready(SimpleBus2AXI4Converter_2_io_in_resp_ready),
    .io_in_resp_valid(SimpleBus2AXI4Converter_2_io_in_resp_valid),
    .io_in_resp_bits_rdata(SimpleBus2AXI4Converter_2_io_in_resp_bits_rdata),
    .io_out_aw_ready(SimpleBus2AXI4Converter_2_io_out_aw_ready),
    .io_out_aw_valid(SimpleBus2AXI4Converter_2_io_out_aw_valid),
    .io_out_aw_bits_addr(SimpleBus2AXI4Converter_2_io_out_aw_bits_addr),
    .io_out_w_ready(SimpleBus2AXI4Converter_2_io_out_w_ready),
    .io_out_w_valid(SimpleBus2AXI4Converter_2_io_out_w_valid),
    .io_out_w_bits_data(SimpleBus2AXI4Converter_2_io_out_w_bits_data),
    .io_out_w_bits_strb(SimpleBus2AXI4Converter_2_io_out_w_bits_strb),
    .io_out_b_ready(SimpleBus2AXI4Converter_2_io_out_b_ready),
    .io_out_b_valid(SimpleBus2AXI4Converter_2_io_out_b_valid),
    .io_out_ar_ready(SimpleBus2AXI4Converter_2_io_out_ar_ready),
    .io_out_ar_valid(SimpleBus2AXI4Converter_2_io_out_ar_valid),
    .io_out_ar_bits_addr(SimpleBus2AXI4Converter_2_io_out_ar_bits_addr),
    .io_out_r_ready(SimpleBus2AXI4Converter_2_io_out_r_ready),
    .io_out_r_valid(SimpleBus2AXI4Converter_2_io_out_r_valid),
    .io_out_r_bits_data(SimpleBus2AXI4Converter_2_io_out_r_bits_data)
  );
  SimpleBus2AXI4Converter_1 SimpleBus2AXI4Converter_3 ( // @[ToAXI4.scala 204:24]
    .clock(SimpleBus2AXI4Converter_3_clock),
    .reset(SimpleBus2AXI4Converter_3_reset),
    .io_in_req_ready(SimpleBus2AXI4Converter_3_io_in_req_ready),
    .io_in_req_valid(SimpleBus2AXI4Converter_3_io_in_req_valid),
    .io_in_req_bits_addr(SimpleBus2AXI4Converter_3_io_in_req_bits_addr),
    .io_in_req_bits_cmd(SimpleBus2AXI4Converter_3_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(SimpleBus2AXI4Converter_3_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(SimpleBus2AXI4Converter_3_io_in_req_bits_wdata),
    .io_in_resp_ready(SimpleBus2AXI4Converter_3_io_in_resp_ready),
    .io_in_resp_valid(SimpleBus2AXI4Converter_3_io_in_resp_valid),
    .io_in_resp_bits_rdata(SimpleBus2AXI4Converter_3_io_in_resp_bits_rdata),
    .io_out_aw_ready(SimpleBus2AXI4Converter_3_io_out_aw_ready),
    .io_out_aw_valid(SimpleBus2AXI4Converter_3_io_out_aw_valid),
    .io_out_aw_bits_addr(SimpleBus2AXI4Converter_3_io_out_aw_bits_addr),
    .io_out_w_ready(SimpleBus2AXI4Converter_3_io_out_w_ready),
    .io_out_w_valid(SimpleBus2AXI4Converter_3_io_out_w_valid),
    .io_out_w_bits_data(SimpleBus2AXI4Converter_3_io_out_w_bits_data),
    .io_out_w_bits_strb(SimpleBus2AXI4Converter_3_io_out_w_bits_strb),
    .io_out_b_ready(SimpleBus2AXI4Converter_3_io_out_b_ready),
    .io_out_b_valid(SimpleBus2AXI4Converter_3_io_out_b_valid),
    .io_out_ar_ready(SimpleBus2AXI4Converter_3_io_out_ar_ready),
    .io_out_ar_valid(SimpleBus2AXI4Converter_3_io_out_ar_valid),
    .io_out_ar_bits_addr(SimpleBus2AXI4Converter_3_io_out_ar_bits_addr),
    .io_out_r_ready(SimpleBus2AXI4Converter_3_io_out_r_ready),
    .io_out_r_valid(SimpleBus2AXI4Converter_3_io_out_r_valid),
    .io_out_r_bits_data(SimpleBus2AXI4Converter_3_io_out_r_bits_data)
  );
  SimpleBus2AXI4Converter_1 SimpleBus2AXI4Converter_4 ( // @[ToAXI4.scala 204:24]
    .clock(SimpleBus2AXI4Converter_4_clock),
    .reset(SimpleBus2AXI4Converter_4_reset),
    .io_in_req_ready(SimpleBus2AXI4Converter_4_io_in_req_ready),
    .io_in_req_valid(SimpleBus2AXI4Converter_4_io_in_req_valid),
    .io_in_req_bits_addr(SimpleBus2AXI4Converter_4_io_in_req_bits_addr),
    .io_in_req_bits_cmd(SimpleBus2AXI4Converter_4_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(SimpleBus2AXI4Converter_4_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(SimpleBus2AXI4Converter_4_io_in_req_bits_wdata),
    .io_in_resp_ready(SimpleBus2AXI4Converter_4_io_in_resp_ready),
    .io_in_resp_valid(SimpleBus2AXI4Converter_4_io_in_resp_valid),
    .io_in_resp_bits_rdata(SimpleBus2AXI4Converter_4_io_in_resp_bits_rdata),
    .io_out_aw_ready(SimpleBus2AXI4Converter_4_io_out_aw_ready),
    .io_out_aw_valid(SimpleBus2AXI4Converter_4_io_out_aw_valid),
    .io_out_aw_bits_addr(SimpleBus2AXI4Converter_4_io_out_aw_bits_addr),
    .io_out_w_ready(SimpleBus2AXI4Converter_4_io_out_w_ready),
    .io_out_w_valid(SimpleBus2AXI4Converter_4_io_out_w_valid),
    .io_out_w_bits_data(SimpleBus2AXI4Converter_4_io_out_w_bits_data),
    .io_out_w_bits_strb(SimpleBus2AXI4Converter_4_io_out_w_bits_strb),
    .io_out_b_ready(SimpleBus2AXI4Converter_4_io_out_b_ready),
    .io_out_b_valid(SimpleBus2AXI4Converter_4_io_out_b_valid),
    .io_out_ar_ready(SimpleBus2AXI4Converter_4_io_out_ar_ready),
    .io_out_ar_valid(SimpleBus2AXI4Converter_4_io_out_ar_valid),
    .io_out_ar_bits_addr(SimpleBus2AXI4Converter_4_io_out_ar_bits_addr),
    .io_out_r_ready(SimpleBus2AXI4Converter_4_io_out_r_ready),
    .io_out_r_valid(SimpleBus2AXI4Converter_4_io_out_r_valid),
    .io_out_r_bits_data(SimpleBus2AXI4Converter_4_io_out_r_bits_data)
  );
  SimpleBus2AXI4Converter_1 SimpleBus2AXI4Converter_5 ( // @[ToAXI4.scala 204:24]
    .clock(SimpleBus2AXI4Converter_5_clock),
    .reset(SimpleBus2AXI4Converter_5_reset),
    .io_in_req_ready(SimpleBus2AXI4Converter_5_io_in_req_ready),
    .io_in_req_valid(SimpleBus2AXI4Converter_5_io_in_req_valid),
    .io_in_req_bits_addr(SimpleBus2AXI4Converter_5_io_in_req_bits_addr),
    .io_in_req_bits_cmd(SimpleBus2AXI4Converter_5_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(SimpleBus2AXI4Converter_5_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(SimpleBus2AXI4Converter_5_io_in_req_bits_wdata),
    .io_in_resp_ready(SimpleBus2AXI4Converter_5_io_in_resp_ready),
    .io_in_resp_valid(SimpleBus2AXI4Converter_5_io_in_resp_valid),
    .io_in_resp_bits_rdata(SimpleBus2AXI4Converter_5_io_in_resp_bits_rdata),
    .io_out_aw_ready(SimpleBus2AXI4Converter_5_io_out_aw_ready),
    .io_out_aw_valid(SimpleBus2AXI4Converter_5_io_out_aw_valid),
    .io_out_aw_bits_addr(SimpleBus2AXI4Converter_5_io_out_aw_bits_addr),
    .io_out_w_ready(SimpleBus2AXI4Converter_5_io_out_w_ready),
    .io_out_w_valid(SimpleBus2AXI4Converter_5_io_out_w_valid),
    .io_out_w_bits_data(SimpleBus2AXI4Converter_5_io_out_w_bits_data),
    .io_out_w_bits_strb(SimpleBus2AXI4Converter_5_io_out_w_bits_strb),
    .io_out_b_ready(SimpleBus2AXI4Converter_5_io_out_b_ready),
    .io_out_b_valid(SimpleBus2AXI4Converter_5_io_out_b_valid),
    .io_out_ar_ready(SimpleBus2AXI4Converter_5_io_out_ar_ready),
    .io_out_ar_valid(SimpleBus2AXI4Converter_5_io_out_ar_valid),
    .io_out_ar_bits_addr(SimpleBus2AXI4Converter_5_io_out_ar_bits_addr),
    .io_out_r_ready(SimpleBus2AXI4Converter_5_io_out_r_ready),
    .io_out_r_valid(SimpleBus2AXI4Converter_5_io_out_r_valid),
    .io_out_r_bits_data(SimpleBus2AXI4Converter_5_io_out_r_bits_data)
  );
  SimpleBus2AXI4Converter_1 SimpleBus2AXI4Converter_6 ( // @[ToAXI4.scala 204:24]
    .clock(SimpleBus2AXI4Converter_6_clock),
    .reset(SimpleBus2AXI4Converter_6_reset),
    .io_in_req_ready(SimpleBus2AXI4Converter_6_io_in_req_ready),
    .io_in_req_valid(SimpleBus2AXI4Converter_6_io_in_req_valid),
    .io_in_req_bits_addr(SimpleBus2AXI4Converter_6_io_in_req_bits_addr),
    .io_in_req_bits_cmd(SimpleBus2AXI4Converter_6_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(SimpleBus2AXI4Converter_6_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(SimpleBus2AXI4Converter_6_io_in_req_bits_wdata),
    .io_in_resp_ready(SimpleBus2AXI4Converter_6_io_in_resp_ready),
    .io_in_resp_valid(SimpleBus2AXI4Converter_6_io_in_resp_valid),
    .io_in_resp_bits_rdata(SimpleBus2AXI4Converter_6_io_in_resp_bits_rdata),
    .io_out_aw_ready(SimpleBus2AXI4Converter_6_io_out_aw_ready),
    .io_out_aw_valid(SimpleBus2AXI4Converter_6_io_out_aw_valid),
    .io_out_aw_bits_addr(SimpleBus2AXI4Converter_6_io_out_aw_bits_addr),
    .io_out_w_ready(SimpleBus2AXI4Converter_6_io_out_w_ready),
    .io_out_w_valid(SimpleBus2AXI4Converter_6_io_out_w_valid),
    .io_out_w_bits_data(SimpleBus2AXI4Converter_6_io_out_w_bits_data),
    .io_out_w_bits_strb(SimpleBus2AXI4Converter_6_io_out_w_bits_strb),
    .io_out_b_ready(SimpleBus2AXI4Converter_6_io_out_b_ready),
    .io_out_b_valid(SimpleBus2AXI4Converter_6_io_out_b_valid),
    .io_out_ar_ready(SimpleBus2AXI4Converter_6_io_out_ar_ready),
    .io_out_ar_valid(SimpleBus2AXI4Converter_6_io_out_ar_valid),
    .io_out_ar_bits_addr(SimpleBus2AXI4Converter_6_io_out_ar_bits_addr),
    .io_out_r_ready(SimpleBus2AXI4Converter_6_io_out_r_ready),
    .io_out_r_valid(SimpleBus2AXI4Converter_6_io_out_r_valid),
    .io_out_r_bits_data(SimpleBus2AXI4Converter_6_io_out_r_bits_data)
  );
  SimpleBus2AXI4Converter_1 SimpleBus2AXI4Converter_7 ( // @[ToAXI4.scala 204:24]
    .clock(SimpleBus2AXI4Converter_7_clock),
    .reset(SimpleBus2AXI4Converter_7_reset),
    .io_in_req_ready(SimpleBus2AXI4Converter_7_io_in_req_ready),
    .io_in_req_valid(SimpleBus2AXI4Converter_7_io_in_req_valid),
    .io_in_req_bits_addr(SimpleBus2AXI4Converter_7_io_in_req_bits_addr),
    .io_in_req_bits_cmd(SimpleBus2AXI4Converter_7_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(SimpleBus2AXI4Converter_7_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(SimpleBus2AXI4Converter_7_io_in_req_bits_wdata),
    .io_in_resp_ready(SimpleBus2AXI4Converter_7_io_in_resp_ready),
    .io_in_resp_valid(SimpleBus2AXI4Converter_7_io_in_resp_valid),
    .io_in_resp_bits_rdata(SimpleBus2AXI4Converter_7_io_in_resp_bits_rdata),
    .io_out_aw_ready(SimpleBus2AXI4Converter_7_io_out_aw_ready),
    .io_out_aw_valid(SimpleBus2AXI4Converter_7_io_out_aw_valid),
    .io_out_aw_bits_addr(SimpleBus2AXI4Converter_7_io_out_aw_bits_addr),
    .io_out_w_ready(SimpleBus2AXI4Converter_7_io_out_w_ready),
    .io_out_w_valid(SimpleBus2AXI4Converter_7_io_out_w_valid),
    .io_out_w_bits_data(SimpleBus2AXI4Converter_7_io_out_w_bits_data),
    .io_out_w_bits_strb(SimpleBus2AXI4Converter_7_io_out_w_bits_strb),
    .io_out_b_ready(SimpleBus2AXI4Converter_7_io_out_b_ready),
    .io_out_b_valid(SimpleBus2AXI4Converter_7_io_out_b_valid),
    .io_out_ar_ready(SimpleBus2AXI4Converter_7_io_out_ar_ready),
    .io_out_ar_valid(SimpleBus2AXI4Converter_7_io_out_ar_valid),
    .io_out_ar_bits_addr(SimpleBus2AXI4Converter_7_io_out_ar_bits_addr),
    .io_out_r_ready(SimpleBus2AXI4Converter_7_io_out_r_ready),
    .io_out_r_valid(SimpleBus2AXI4Converter_7_io_out_r_valid),
    .io_out_r_bits_data(SimpleBus2AXI4Converter_7_io_out_r_bits_data)
  );
  assign io_rw_req_ready = xbar_io_in_req_ready; // @[SimMMIO.scala 46:14]
  assign io_rw_resp_valid = xbar_io_in_resp_valid; // @[SimMMIO.scala 46:14]
  assign io_rw_resp_bits_rdata = xbar_io_in_resp_bits_rdata; // @[SimMMIO.scala 46:14]
  assign io_difftestCtrl_enable = difftestCtrl_io_extra_enable; // @[SimMMIO.scala 64:19]
  assign io_meip = meipGen_io_extra_enable; // @[SimMMIO.scala 65:11]
  assign io_dma_aw_valid = dma_io_extra_dma_aw_valid; // @[SimMMIO.scala 63:10]
  assign io_dma_aw_bits_addr = dma_io_extra_dma_aw_bits_addr; // @[SimMMIO.scala 63:10]
  assign io_dma_aw_bits_len = dma_io_extra_dma_aw_bits_len; // @[SimMMIO.scala 63:10]
  assign io_dma_aw_bits_size = dma_io_extra_dma_aw_bits_size; // @[SimMMIO.scala 63:10]
  assign io_dma_w_valid = dma_io_extra_dma_w_valid; // @[SimMMIO.scala 63:10]
  assign io_dma_w_bits_data = dma_io_extra_dma_w_bits_data; // @[SimMMIO.scala 63:10]
  assign io_dma_w_bits_strb = dma_io_extra_dma_w_bits_strb; // @[SimMMIO.scala 63:10]
  assign io_dma_b_ready = dma_io_extra_dma_b_ready; // @[SimMMIO.scala 63:10]
  assign io_dma_ar_valid = dma_io_extra_dma_ar_valid; // @[SimMMIO.scala 63:10]
  assign io_dma_ar_bits_addr = dma_io_extra_dma_ar_bits_addr; // @[SimMMIO.scala 63:10]
  assign io_dma_r_ready = dma_io_extra_dma_r_ready; // @[SimMMIO.scala 63:10]
  assign xbar_clock = clock;
  assign xbar_reset = reset;
  assign xbar_io_in_req_valid = io_rw_req_valid; // @[SimMMIO.scala 46:14]
  assign xbar_io_in_req_bits_addr = io_rw_req_bits_addr; // @[SimMMIO.scala 46:14]
  assign xbar_io_in_req_bits_size = io_rw_req_bits_size; // @[SimMMIO.scala 46:14]
  assign xbar_io_in_req_bits_cmd = io_rw_req_bits_cmd; // @[SimMMIO.scala 46:14]
  assign xbar_io_in_req_bits_wmask = io_rw_req_bits_wmask; // @[SimMMIO.scala 46:14]
  assign xbar_io_in_req_bits_wdata = io_rw_req_bits_wdata; // @[SimMMIO.scala 46:14]
  assign xbar_io_in_resp_ready = io_rw_resp_ready; // @[SimMMIO.scala 46:14]
  assign xbar_io_out_0_req_ready = SimpleBus2AXI4Converter_io_in_req_ready; // @[ToAXI4.scala 205:18]
  assign xbar_io_out_0_resp_valid = SimpleBus2AXI4Converter_io_in_resp_valid; // @[ToAXI4.scala 205:18]
  assign xbar_io_out_0_resp_bits_rdata = SimpleBus2AXI4Converter_io_in_resp_bits_rdata; // @[ToAXI4.scala 205:18]
  assign xbar_io_out_1_req_ready = SimpleBus2AXI4Converter_1_io_in_req_ready; // @[ToAXI4.scala 205:18]
  assign xbar_io_out_1_resp_valid = SimpleBus2AXI4Converter_1_io_in_resp_valid; // @[ToAXI4.scala 205:18]
  assign xbar_io_out_1_resp_bits_rdata = SimpleBus2AXI4Converter_1_io_in_resp_bits_rdata; // @[ToAXI4.scala 205:18]
  assign xbar_io_out_2_req_ready = SimpleBus2AXI4Converter_2_io_in_req_ready; // @[ToAXI4.scala 205:18]
  assign xbar_io_out_2_resp_valid = SimpleBus2AXI4Converter_2_io_in_resp_valid; // @[ToAXI4.scala 205:18]
  assign xbar_io_out_2_resp_bits_rdata = SimpleBus2AXI4Converter_2_io_in_resp_bits_rdata; // @[ToAXI4.scala 205:18]
  assign xbar_io_out_3_req_ready = SimpleBus2AXI4Converter_3_io_in_req_ready; // @[ToAXI4.scala 205:18]
  assign xbar_io_out_3_resp_valid = SimpleBus2AXI4Converter_3_io_in_resp_valid; // @[ToAXI4.scala 205:18]
  assign xbar_io_out_3_resp_bits_rdata = SimpleBus2AXI4Converter_3_io_in_resp_bits_rdata; // @[ToAXI4.scala 205:18]
  assign xbar_io_out_4_req_ready = SimpleBus2AXI4Converter_4_io_in_req_ready; // @[ToAXI4.scala 205:18]
  assign xbar_io_out_4_resp_valid = SimpleBus2AXI4Converter_4_io_in_resp_valid; // @[ToAXI4.scala 205:18]
  assign xbar_io_out_4_resp_bits_rdata = SimpleBus2AXI4Converter_4_io_in_resp_bits_rdata; // @[ToAXI4.scala 205:18]
  assign xbar_io_out_5_req_ready = SimpleBus2AXI4Converter_5_io_in_req_ready; // @[ToAXI4.scala 205:18]
  assign xbar_io_out_5_resp_valid = SimpleBus2AXI4Converter_5_io_in_resp_valid; // @[ToAXI4.scala 205:18]
  assign xbar_io_out_5_resp_bits_rdata = SimpleBus2AXI4Converter_5_io_in_resp_bits_rdata; // @[ToAXI4.scala 205:18]
  assign xbar_io_out_6_req_ready = SimpleBus2AXI4Converter_6_io_in_req_ready; // @[ToAXI4.scala 205:18]
  assign xbar_io_out_6_resp_valid = SimpleBus2AXI4Converter_6_io_in_resp_valid; // @[ToAXI4.scala 205:18]
  assign xbar_io_out_6_resp_bits_rdata = SimpleBus2AXI4Converter_6_io_in_resp_bits_rdata; // @[ToAXI4.scala 205:18]
  assign xbar_io_out_7_req_ready = SimpleBus2AXI4Converter_7_io_in_req_ready; // @[ToAXI4.scala 205:18]
  assign xbar_io_out_7_resp_valid = SimpleBus2AXI4Converter_7_io_in_resp_valid; // @[ToAXI4.scala 205:18]
  assign xbar_io_out_7_resp_bits_rdata = SimpleBus2AXI4Converter_7_io_in_resp_bits_rdata; // @[ToAXI4.scala 205:18]
  assign xbar_DISPLAY_ENABLE = _T_13;
  assign uart_clock = clock;
  assign uart_reset = reset;
  assign uart_io_in_aw_valid = SimpleBus2AXI4Converter_io_out_aw_valid; // @[SimMMIO.scala 55:14]
  assign uart_io_in_aw_bits_addr = SimpleBus2AXI4Converter_io_out_aw_bits_addr; // @[SimMMIO.scala 55:14]
  assign uart_io_in_w_valid = SimpleBus2AXI4Converter_io_out_w_valid; // @[SimMMIO.scala 55:14]
  assign uart_io_in_w_bits_data = SimpleBus2AXI4Converter_io_out_w_bits_data; // @[SimMMIO.scala 55:14]
  assign uart_io_in_w_bits_strb = SimpleBus2AXI4Converter_io_out_w_bits_strb; // @[SimMMIO.scala 55:14]
  assign uart_io_in_b_ready = SimpleBus2AXI4Converter_io_out_b_ready; // @[SimMMIO.scala 55:14]
  assign uart_io_in_ar_valid = SimpleBus2AXI4Converter_io_out_ar_valid; // @[SimMMIO.scala 55:14]
  assign uart_io_in_ar_bits_addr = SimpleBus2AXI4Converter_io_out_ar_bits_addr; // @[SimMMIO.scala 55:14]
  assign uart_io_in_r_ready = SimpleBus2AXI4Converter_io_out_r_ready; // @[SimMMIO.scala 55:14]
  assign vga_clock = clock;
  assign vga_reset = reset;
  assign vga_io_in_fb_aw_valid = SimpleBus2AXI4Converter_1_io_out_aw_valid; // @[SimMMIO.scala 56:16]
  assign vga_io_in_fb_aw_bits_addr = SimpleBus2AXI4Converter_1_io_out_aw_bits_addr; // @[SimMMIO.scala 56:16]
  assign vga_io_in_fb_w_valid = SimpleBus2AXI4Converter_1_io_out_w_valid; // @[SimMMIO.scala 56:16]
  assign vga_io_in_fb_w_bits_data = SimpleBus2AXI4Converter_1_io_out_w_bits_data; // @[SimMMIO.scala 56:16]
  assign vga_io_in_fb_w_bits_strb = SimpleBus2AXI4Converter_1_io_out_w_bits_strb; // @[SimMMIO.scala 56:16]
  assign vga_io_in_fb_b_ready = SimpleBus2AXI4Converter_1_io_out_b_ready; // @[SimMMIO.scala 56:16]
  assign vga_io_in_fb_ar_valid = SimpleBus2AXI4Converter_1_io_out_ar_valid; // @[SimMMIO.scala 56:16]
  assign vga_io_in_fb_r_ready = SimpleBus2AXI4Converter_1_io_out_r_ready; // @[SimMMIO.scala 56:16]
  assign vga_io_in_ctrl_aw_valid = SimpleBus2AXI4Converter_2_io_out_aw_valid; // @[SimMMIO.scala 57:18]
  assign vga_io_in_ctrl_w_valid = SimpleBus2AXI4Converter_2_io_out_w_valid; // @[SimMMIO.scala 57:18]
  assign vga_io_in_ctrl_b_ready = SimpleBus2AXI4Converter_2_io_out_b_ready; // @[SimMMIO.scala 57:18]
  assign vga_io_in_ctrl_ar_valid = SimpleBus2AXI4Converter_2_io_out_ar_valid; // @[SimMMIO.scala 57:18]
  assign vga_io_in_ctrl_ar_bits_addr = SimpleBus2AXI4Converter_2_io_out_ar_bits_addr; // @[SimMMIO.scala 57:18]
  assign vga_io_in_ctrl_r_ready = SimpleBus2AXI4Converter_2_io_out_r_ready; // @[SimMMIO.scala 57:18]
  assign flash_clock = clock;
  assign flash_reset = reset;
  assign flash_io_in_aw_valid = SimpleBus2AXI4Converter_3_io_out_aw_valid; // @[SimMMIO.scala 58:15]
  assign flash_io_in_w_valid = SimpleBus2AXI4Converter_3_io_out_w_valid; // @[SimMMIO.scala 58:15]
  assign flash_io_in_b_ready = SimpleBus2AXI4Converter_3_io_out_b_ready; // @[SimMMIO.scala 58:15]
  assign flash_io_in_ar_valid = SimpleBus2AXI4Converter_3_io_out_ar_valid; // @[SimMMIO.scala 58:15]
  assign flash_io_in_ar_bits_addr = SimpleBus2AXI4Converter_3_io_out_ar_bits_addr; // @[SimMMIO.scala 58:15]
  assign flash_io_in_r_ready = SimpleBus2AXI4Converter_3_io_out_r_ready; // @[SimMMIO.scala 58:15]
  assign sd_clock = clock;
  assign sd_reset = reset;
  assign sd_io_in_aw_valid = SimpleBus2AXI4Converter_4_io_out_aw_valid; // @[SimMMIO.scala 59:12]
  assign sd_io_in_aw_bits_addr = SimpleBus2AXI4Converter_4_io_out_aw_bits_addr; // @[SimMMIO.scala 59:12]
  assign sd_io_in_w_valid = SimpleBus2AXI4Converter_4_io_out_w_valid; // @[SimMMIO.scala 59:12]
  assign sd_io_in_w_bits_data = SimpleBus2AXI4Converter_4_io_out_w_bits_data; // @[SimMMIO.scala 59:12]
  assign sd_io_in_w_bits_strb = SimpleBus2AXI4Converter_4_io_out_w_bits_strb; // @[SimMMIO.scala 59:12]
  assign sd_io_in_b_ready = SimpleBus2AXI4Converter_4_io_out_b_ready; // @[SimMMIO.scala 59:12]
  assign sd_io_in_ar_valid = SimpleBus2AXI4Converter_4_io_out_ar_valid; // @[SimMMIO.scala 59:12]
  assign sd_io_in_ar_bits_addr = SimpleBus2AXI4Converter_4_io_out_ar_bits_addr; // @[SimMMIO.scala 59:12]
  assign sd_io_in_r_ready = SimpleBus2AXI4Converter_4_io_out_r_ready; // @[SimMMIO.scala 59:12]
  assign difftestCtrl_clock = clock;
  assign difftestCtrl_reset = reset;
  assign difftestCtrl_io_in_aw_valid = SimpleBus2AXI4Converter_5_io_out_aw_valid; // @[SimMMIO.scala 60:22]
  assign difftestCtrl_io_in_aw_bits_addr = SimpleBus2AXI4Converter_5_io_out_aw_bits_addr; // @[SimMMIO.scala 60:22]
  assign difftestCtrl_io_in_w_valid = SimpleBus2AXI4Converter_5_io_out_w_valid; // @[SimMMIO.scala 60:22]
  assign difftestCtrl_io_in_w_bits_data = SimpleBus2AXI4Converter_5_io_out_w_bits_data; // @[SimMMIO.scala 60:22]
  assign difftestCtrl_io_in_w_bits_strb = SimpleBus2AXI4Converter_5_io_out_w_bits_strb; // @[SimMMIO.scala 60:22]
  assign difftestCtrl_io_in_b_ready = SimpleBus2AXI4Converter_5_io_out_b_ready; // @[SimMMIO.scala 60:22]
  assign difftestCtrl_io_in_ar_valid = SimpleBus2AXI4Converter_5_io_out_ar_valid; // @[SimMMIO.scala 60:22]
  assign difftestCtrl_io_in_r_ready = SimpleBus2AXI4Converter_5_io_out_r_ready; // @[SimMMIO.scala 60:22]
  assign meipGen_clock = clock;
  assign meipGen_reset = reset;
  assign meipGen_io_in_aw_valid = SimpleBus2AXI4Converter_6_io_out_aw_valid; // @[SimMMIO.scala 61:17]
  assign meipGen_io_in_aw_bits_addr = SimpleBus2AXI4Converter_6_io_out_aw_bits_addr; // @[SimMMIO.scala 61:17]
  assign meipGen_io_in_w_valid = SimpleBus2AXI4Converter_6_io_out_w_valid; // @[SimMMIO.scala 61:17]
  assign meipGen_io_in_w_bits_data = SimpleBus2AXI4Converter_6_io_out_w_bits_data; // @[SimMMIO.scala 61:17]
  assign meipGen_io_in_w_bits_strb = SimpleBus2AXI4Converter_6_io_out_w_bits_strb; // @[SimMMIO.scala 61:17]
  assign meipGen_io_in_b_ready = SimpleBus2AXI4Converter_6_io_out_b_ready; // @[SimMMIO.scala 61:17]
  assign meipGen_io_in_ar_valid = SimpleBus2AXI4Converter_6_io_out_ar_valid; // @[SimMMIO.scala 61:17]
  assign meipGen_io_in_r_ready = SimpleBus2AXI4Converter_6_io_out_r_ready; // @[SimMMIO.scala 61:17]
  assign dma_clock = clock;
  assign dma_reset = reset;
  assign dma_io_in_aw_valid = SimpleBus2AXI4Converter_7_io_out_aw_valid; // @[SimMMIO.scala 62:13]
  assign dma_io_in_aw_bits_addr = SimpleBus2AXI4Converter_7_io_out_aw_bits_addr; // @[SimMMIO.scala 62:13]
  assign dma_io_in_w_valid = SimpleBus2AXI4Converter_7_io_out_w_valid; // @[SimMMIO.scala 62:13]
  assign dma_io_in_w_bits_data = SimpleBus2AXI4Converter_7_io_out_w_bits_data; // @[SimMMIO.scala 62:13]
  assign dma_io_in_w_bits_strb = SimpleBus2AXI4Converter_7_io_out_w_bits_strb; // @[SimMMIO.scala 62:13]
  assign dma_io_in_b_ready = SimpleBus2AXI4Converter_7_io_out_b_ready; // @[SimMMIO.scala 62:13]
  assign dma_io_in_ar_valid = SimpleBus2AXI4Converter_7_io_out_ar_valid; // @[SimMMIO.scala 62:13]
  assign dma_io_in_ar_bits_addr = SimpleBus2AXI4Converter_7_io_out_ar_bits_addr; // @[SimMMIO.scala 62:13]
  assign dma_io_in_r_ready = SimpleBus2AXI4Converter_7_io_out_r_ready; // @[SimMMIO.scala 62:13]
  assign dma_io_extra_dma_aw_ready = io_dma_aw_ready; // @[SimMMIO.scala 63:10]
  assign dma_io_extra_dma_w_ready = io_dma_w_ready; // @[SimMMIO.scala 63:10]
  assign dma_io_extra_dma_b_valid = io_dma_b_valid; // @[SimMMIO.scala 63:10]
  assign dma_io_extra_dma_ar_ready = io_dma_ar_ready; // @[SimMMIO.scala 63:10]
  assign dma_io_extra_dma_r_valid = io_dma_r_valid; // @[SimMMIO.scala 63:10]
  assign dma_io_extra_dma_r_bits_data = io_dma_r_bits_data; // @[SimMMIO.scala 63:10]
  assign SimpleBus2AXI4Converter_clock = clock;
  assign SimpleBus2AXI4Converter_reset = reset;
  assign SimpleBus2AXI4Converter_io_in_req_valid = xbar_io_out_0_req_valid; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_io_in_req_bits_addr = xbar_io_out_0_req_bits_addr; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_io_in_req_bits_cmd = xbar_io_out_0_req_bits_cmd; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_io_in_req_bits_wmask = xbar_io_out_0_req_bits_wmask; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_io_in_req_bits_wdata = xbar_io_out_0_req_bits_wdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_io_in_resp_ready = xbar_io_out_0_resp_ready; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_io_out_aw_ready = uart_io_in_aw_ready; // @[SimMMIO.scala 55:14]
  assign SimpleBus2AXI4Converter_io_out_w_ready = uart_io_in_w_ready; // @[SimMMIO.scala 55:14]
  assign SimpleBus2AXI4Converter_io_out_b_valid = uart_io_in_b_valid; // @[SimMMIO.scala 55:14]
  assign SimpleBus2AXI4Converter_io_out_ar_ready = uart_io_in_ar_ready; // @[SimMMIO.scala 55:14]
  assign SimpleBus2AXI4Converter_io_out_r_valid = uart_io_in_r_valid; // @[SimMMIO.scala 55:14]
  assign SimpleBus2AXI4Converter_io_out_r_bits_data = uart_io_in_r_bits_data; // @[SimMMIO.scala 55:14]
  assign SimpleBus2AXI4Converter_1_clock = clock;
  assign SimpleBus2AXI4Converter_1_reset = reset;
  assign SimpleBus2AXI4Converter_1_io_in_req_valid = xbar_io_out_1_req_valid; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_req_bits_addr = xbar_io_out_1_req_bits_addr; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_req_bits_cmd = xbar_io_out_1_req_bits_cmd; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_req_bits_wmask = xbar_io_out_1_req_bits_wmask; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_req_bits_wdata = xbar_io_out_1_req_bits_wdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_resp_ready = xbar_io_out_1_resp_ready; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_out_aw_ready = vga_io_in_fb_aw_ready; // @[SimMMIO.scala 56:16]
  assign SimpleBus2AXI4Converter_1_io_out_w_ready = vga_io_in_fb_w_ready; // @[SimMMIO.scala 56:16]
  assign SimpleBus2AXI4Converter_1_io_out_b_valid = vga_io_in_fb_b_valid; // @[SimMMIO.scala 56:16]
  assign SimpleBus2AXI4Converter_1_io_out_ar_ready = 1'h1; // @[SimMMIO.scala 56:16]
  assign SimpleBus2AXI4Converter_1_io_out_r_valid = vga_io_in_fb_r_valid; // @[SimMMIO.scala 56:16]
  assign SimpleBus2AXI4Converter_1_io_out_r_bits_data = 64'h0; // @[SimMMIO.scala 56:16]
  assign SimpleBus2AXI4Converter_2_clock = clock;
  assign SimpleBus2AXI4Converter_2_reset = reset;
  assign SimpleBus2AXI4Converter_2_io_in_req_valid = xbar_io_out_2_req_valid; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_in_req_bits_addr = xbar_io_out_2_req_bits_addr; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_in_req_bits_cmd = xbar_io_out_2_req_bits_cmd; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_in_req_bits_wmask = xbar_io_out_2_req_bits_wmask; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_in_req_bits_wdata = xbar_io_out_2_req_bits_wdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_in_resp_ready = xbar_io_out_2_resp_ready; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_out_aw_ready = vga_io_in_ctrl_aw_ready; // @[SimMMIO.scala 57:18]
  assign SimpleBus2AXI4Converter_2_io_out_w_ready = vga_io_in_ctrl_w_ready; // @[SimMMIO.scala 57:18]
  assign SimpleBus2AXI4Converter_2_io_out_b_valid = vga_io_in_ctrl_b_valid; // @[SimMMIO.scala 57:18]
  assign SimpleBus2AXI4Converter_2_io_out_ar_ready = vga_io_in_ctrl_ar_ready; // @[SimMMIO.scala 57:18]
  assign SimpleBus2AXI4Converter_2_io_out_r_valid = vga_io_in_ctrl_r_valid; // @[SimMMIO.scala 57:18]
  assign SimpleBus2AXI4Converter_2_io_out_r_bits_data = vga_io_in_ctrl_r_bits_data; // @[SimMMIO.scala 57:18]
  assign SimpleBus2AXI4Converter_3_clock = clock;
  assign SimpleBus2AXI4Converter_3_reset = reset;
  assign SimpleBus2AXI4Converter_3_io_in_req_valid = xbar_io_out_3_req_valid; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_3_io_in_req_bits_addr = xbar_io_out_3_req_bits_addr; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_3_io_in_req_bits_cmd = xbar_io_out_3_req_bits_cmd; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_3_io_in_req_bits_wmask = xbar_io_out_3_req_bits_wmask; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_3_io_in_req_bits_wdata = xbar_io_out_3_req_bits_wdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_3_io_in_resp_ready = xbar_io_out_3_resp_ready; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_3_io_out_aw_ready = flash_io_in_aw_ready; // @[SimMMIO.scala 58:15]
  assign SimpleBus2AXI4Converter_3_io_out_w_ready = flash_io_in_w_ready; // @[SimMMIO.scala 58:15]
  assign SimpleBus2AXI4Converter_3_io_out_b_valid = flash_io_in_b_valid; // @[SimMMIO.scala 58:15]
  assign SimpleBus2AXI4Converter_3_io_out_ar_ready = flash_io_in_ar_ready; // @[SimMMIO.scala 58:15]
  assign SimpleBus2AXI4Converter_3_io_out_r_valid = flash_io_in_r_valid; // @[SimMMIO.scala 58:15]
  assign SimpleBus2AXI4Converter_3_io_out_r_bits_data = flash_io_in_r_bits_data; // @[SimMMIO.scala 58:15]
  assign SimpleBus2AXI4Converter_4_clock = clock;
  assign SimpleBus2AXI4Converter_4_reset = reset;
  assign SimpleBus2AXI4Converter_4_io_in_req_valid = xbar_io_out_4_req_valid; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_4_io_in_req_bits_addr = xbar_io_out_4_req_bits_addr; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_4_io_in_req_bits_cmd = xbar_io_out_4_req_bits_cmd; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_4_io_in_req_bits_wmask = xbar_io_out_4_req_bits_wmask; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_4_io_in_req_bits_wdata = xbar_io_out_4_req_bits_wdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_4_io_in_resp_ready = xbar_io_out_4_resp_ready; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_4_io_out_aw_ready = sd_io_in_aw_ready; // @[SimMMIO.scala 59:12]
  assign SimpleBus2AXI4Converter_4_io_out_w_ready = sd_io_in_w_ready; // @[SimMMIO.scala 59:12]
  assign SimpleBus2AXI4Converter_4_io_out_b_valid = sd_io_in_b_valid; // @[SimMMIO.scala 59:12]
  assign SimpleBus2AXI4Converter_4_io_out_ar_ready = sd_io_in_ar_ready; // @[SimMMIO.scala 59:12]
  assign SimpleBus2AXI4Converter_4_io_out_r_valid = sd_io_in_r_valid; // @[SimMMIO.scala 59:12]
  assign SimpleBus2AXI4Converter_4_io_out_r_bits_data = sd_io_in_r_bits_data; // @[SimMMIO.scala 59:12]
  assign SimpleBus2AXI4Converter_5_clock = clock;
  assign SimpleBus2AXI4Converter_5_reset = reset;
  assign SimpleBus2AXI4Converter_5_io_in_req_valid = xbar_io_out_5_req_valid; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_5_io_in_req_bits_addr = xbar_io_out_5_req_bits_addr; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_5_io_in_req_bits_cmd = xbar_io_out_5_req_bits_cmd; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_5_io_in_req_bits_wmask = xbar_io_out_5_req_bits_wmask; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_5_io_in_req_bits_wdata = xbar_io_out_5_req_bits_wdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_5_io_in_resp_ready = xbar_io_out_5_resp_ready; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_5_io_out_aw_ready = difftestCtrl_io_in_aw_ready; // @[SimMMIO.scala 60:22]
  assign SimpleBus2AXI4Converter_5_io_out_w_ready = difftestCtrl_io_in_w_ready; // @[SimMMIO.scala 60:22]
  assign SimpleBus2AXI4Converter_5_io_out_b_valid = difftestCtrl_io_in_b_valid; // @[SimMMIO.scala 60:22]
  assign SimpleBus2AXI4Converter_5_io_out_ar_ready = difftestCtrl_io_in_ar_ready; // @[SimMMIO.scala 60:22]
  assign SimpleBus2AXI4Converter_5_io_out_r_valid = difftestCtrl_io_in_r_valid; // @[SimMMIO.scala 60:22]
  assign SimpleBus2AXI4Converter_5_io_out_r_bits_data = difftestCtrl_io_in_r_bits_data; // @[SimMMIO.scala 60:22]
  assign SimpleBus2AXI4Converter_6_clock = clock;
  assign SimpleBus2AXI4Converter_6_reset = reset;
  assign SimpleBus2AXI4Converter_6_io_in_req_valid = xbar_io_out_6_req_valid; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_6_io_in_req_bits_addr = xbar_io_out_6_req_bits_addr; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_6_io_in_req_bits_cmd = xbar_io_out_6_req_bits_cmd; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_6_io_in_req_bits_wmask = xbar_io_out_6_req_bits_wmask; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_6_io_in_req_bits_wdata = xbar_io_out_6_req_bits_wdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_6_io_in_resp_ready = xbar_io_out_6_resp_ready; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_6_io_out_aw_ready = meipGen_io_in_aw_ready; // @[SimMMIO.scala 61:17]
  assign SimpleBus2AXI4Converter_6_io_out_w_ready = meipGen_io_in_w_ready; // @[SimMMIO.scala 61:17]
  assign SimpleBus2AXI4Converter_6_io_out_b_valid = meipGen_io_in_b_valid; // @[SimMMIO.scala 61:17]
  assign SimpleBus2AXI4Converter_6_io_out_ar_ready = meipGen_io_in_ar_ready; // @[SimMMIO.scala 61:17]
  assign SimpleBus2AXI4Converter_6_io_out_r_valid = meipGen_io_in_r_valid; // @[SimMMIO.scala 61:17]
  assign SimpleBus2AXI4Converter_6_io_out_r_bits_data = meipGen_io_in_r_bits_data; // @[SimMMIO.scala 61:17]
  assign SimpleBus2AXI4Converter_7_clock = clock;
  assign SimpleBus2AXI4Converter_7_reset = reset;
  assign SimpleBus2AXI4Converter_7_io_in_req_valid = xbar_io_out_7_req_valid; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_7_io_in_req_bits_addr = xbar_io_out_7_req_bits_addr; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_7_io_in_req_bits_cmd = xbar_io_out_7_req_bits_cmd; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_7_io_in_req_bits_wmask = xbar_io_out_7_req_bits_wmask; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_7_io_in_req_bits_wdata = xbar_io_out_7_req_bits_wdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_7_io_in_resp_ready = xbar_io_out_7_resp_ready; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_7_io_out_aw_ready = dma_io_in_aw_ready; // @[SimMMIO.scala 62:13]
  assign SimpleBus2AXI4Converter_7_io_out_w_ready = dma_io_in_w_ready; // @[SimMMIO.scala 62:13]
  assign SimpleBus2AXI4Converter_7_io_out_b_valid = dma_io_in_b_valid; // @[SimMMIO.scala 62:13]
  assign SimpleBus2AXI4Converter_7_io_out_ar_ready = dma_io_in_ar_ready; // @[SimMMIO.scala 62:13]
  assign SimpleBus2AXI4Converter_7_io_out_r_valid = dma_io_in_r_valid; // @[SimMMIO.scala 62:13]
  assign SimpleBus2AXI4Converter_7_io_out_r_bits_data = dma_io_in_r_bits_data; // @[SimMMIO.scala 62:13]
endmodule
module NutShellSimTop(
  input         clock,
  input         reset,
  output [63:0] io_difftest_r_0,
  output [63:0] io_difftest_r_1,
  output [63:0] io_difftest_r_2,
  output [63:0] io_difftest_r_3,
  output [63:0] io_difftest_r_4,
  output [63:0] io_difftest_r_5,
  output [63:0] io_difftest_r_6,
  output [63:0] io_difftest_r_7,
  output [63:0] io_difftest_r_8,
  output [63:0] io_difftest_r_9,
  output [63:0] io_difftest_r_10,
  output [63:0] io_difftest_r_11,
  output [63:0] io_difftest_r_12,
  output [63:0] io_difftest_r_13,
  output [63:0] io_difftest_r_14,
  output [63:0] io_difftest_r_15,
  output [63:0] io_difftest_r_16,
  output [63:0] io_difftest_r_17,
  output [63:0] io_difftest_r_18,
  output [63:0] io_difftest_r_19,
  output [63:0] io_difftest_r_20,
  output [63:0] io_difftest_r_21,
  output [63:0] io_difftest_r_22,
  output [63:0] io_difftest_r_23,
  output [63:0] io_difftest_r_24,
  output [63:0] io_difftest_r_25,
  output [63:0] io_difftest_r_26,
  output [63:0] io_difftest_r_27,
  output [63:0] io_difftest_r_28,
  output [63:0] io_difftest_r_29,
  output [63:0] io_difftest_r_30,
  output [63:0] io_difftest_r_31,
  output [63:0] io_difftest_sr_0,
  output [63:0] io_difftest_sr_1,
  output [63:0] io_difftest_sr_2,
  output [63:0] io_difftest_sr_3,
  output [63:0] io_difftest_sr_4,
  output        io_difftest_commit,
  output        io_difftest_isMultiCommit,
  output [63:0] io_difftest_thisPC,
  output [31:0] io_difftest_thisINST,
  output        io_difftest_isMMIO,
  output        io_difftest_isRVC,
  output        io_difftest_isRVC2,
  output [63:0] io_difftest_intrNO,
  output [1:0]  io_difftest_priviledgeMode,
  output [63:0] io_difftest_mstatus,
  output [63:0] io_difftest_sstatus,
  output [63:0] io_difftest_mepc,
  output [63:0] io_difftest_sepc,
  output [63:0] io_difftest_mcause,
  output [63:0] io_difftest_scause,
  input  [63:0] io_logCtrl_log_begin,
  input  [63:0] io_logCtrl_log_end,
  input  [63:0] io_logCtrl_log_level,
  output        io_difftestCtrl_enable
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  soc_clock; // @[NutShellSim.scala 65:19]
  wire  soc_reset; // @[NutShellSim.scala 65:19]
  wire  soc_io_mem_aw_ready; // @[NutShellSim.scala 65:19]
  wire  soc_io_mem_aw_valid; // @[NutShellSim.scala 65:19]
  wire [31:0] soc_io_mem_aw_bits_addr; // @[NutShellSim.scala 65:19]
  wire [7:0] soc_io_mem_aw_bits_len; // @[NutShellSim.scala 65:19]
  wire [2:0] soc_io_mem_aw_bits_size; // @[NutShellSim.scala 65:19]
  wire [1:0] soc_io_mem_aw_bits_burst; // @[NutShellSim.scala 65:19]
  wire  soc_io_mem_w_ready; // @[NutShellSim.scala 65:19]
  wire  soc_io_mem_w_valid; // @[NutShellSim.scala 65:19]
  wire [63:0] soc_io_mem_w_bits_data; // @[NutShellSim.scala 65:19]
  wire  soc_io_mem_w_bits_last; // @[NutShellSim.scala 65:19]
  wire  soc_io_mem_b_valid; // @[NutShellSim.scala 65:19]
  wire  soc_io_mem_ar_ready; // @[NutShellSim.scala 65:19]
  wire  soc_io_mem_ar_valid; // @[NutShellSim.scala 65:19]
  wire [31:0] soc_io_mem_ar_bits_addr; // @[NutShellSim.scala 65:19]
  wire [7:0] soc_io_mem_ar_bits_len; // @[NutShellSim.scala 65:19]
  wire  soc_io_mem_r_valid; // @[NutShellSim.scala 65:19]
  wire [63:0] soc_io_mem_r_bits_data; // @[NutShellSim.scala 65:19]
  wire  soc_io_mem_r_bits_last; // @[NutShellSim.scala 65:19]
  wire  soc_io_mmio_req_ready; // @[NutShellSim.scala 65:19]
  wire  soc_io_mmio_req_valid; // @[NutShellSim.scala 65:19]
  wire [31:0] soc_io_mmio_req_bits_addr; // @[NutShellSim.scala 65:19]
  wire [2:0] soc_io_mmio_req_bits_size; // @[NutShellSim.scala 65:19]
  wire [3:0] soc_io_mmio_req_bits_cmd; // @[NutShellSim.scala 65:19]
  wire [7:0] soc_io_mmio_req_bits_wmask; // @[NutShellSim.scala 65:19]
  wire [63:0] soc_io_mmio_req_bits_wdata; // @[NutShellSim.scala 65:19]
  wire  soc_io_mmio_resp_ready; // @[NutShellSim.scala 65:19]
  wire  soc_io_mmio_resp_valid; // @[NutShellSim.scala 65:19]
  wire [63:0] soc_io_mmio_resp_bits_rdata; // @[NutShellSim.scala 65:19]
  wire  soc_io_frontend_aw_ready; // @[NutShellSim.scala 65:19]
  wire  soc_io_frontend_aw_valid; // @[NutShellSim.scala 65:19]
  wire [31:0] soc_io_frontend_aw_bits_addr; // @[NutShellSim.scala 65:19]
  wire [7:0] soc_io_frontend_aw_bits_len; // @[NutShellSim.scala 65:19]
  wire [2:0] soc_io_frontend_aw_bits_size; // @[NutShellSim.scala 65:19]
  wire  soc_io_frontend_w_ready; // @[NutShellSim.scala 65:19]
  wire  soc_io_frontend_w_valid; // @[NutShellSim.scala 65:19]
  wire [63:0] soc_io_frontend_w_bits_data; // @[NutShellSim.scala 65:19]
  wire [7:0] soc_io_frontend_w_bits_strb; // @[NutShellSim.scala 65:19]
  wire  soc_io_frontend_b_ready; // @[NutShellSim.scala 65:19]
  wire  soc_io_frontend_b_valid; // @[NutShellSim.scala 65:19]
  wire  soc_io_frontend_ar_ready; // @[NutShellSim.scala 65:19]
  wire  soc_io_frontend_ar_valid; // @[NutShellSim.scala 65:19]
  wire [31:0] soc_io_frontend_ar_bits_addr; // @[NutShellSim.scala 65:19]
  wire  soc_io_frontend_r_ready; // @[NutShellSim.scala 65:19]
  wire  soc_io_frontend_r_valid; // @[NutShellSim.scala 65:19]
  wire [63:0] soc_io_frontend_r_bits_data; // @[NutShellSim.scala 65:19]
  wire  soc_io_meip; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_4181; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_4184; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_4185; // @[NutShellSim.scala 65:19]
  wire  soc_falseWire; // @[NutShellSim.scala 65:19]
  wire  soc_falseWire_0; // @[NutShellSim.scala 65:19]
  wire [1:0] soc__T_4178; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_284_0; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_284_1; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_284_2; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_284_3; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_284_4; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_284_5; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_284_6; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_284_7; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_284_8; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_284_9; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_284_10; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_284_11; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_284_12; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_284_13; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_284_14; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_284_15; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_284_16; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_284_17; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_284_18; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_284_19; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_284_20; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_284_21; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_284_22; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_284_23; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_284_24; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_284_25; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_284_26; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_284_27; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_284_28; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_284_29; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_284_30; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_284_31; // @[NutShellSim.scala 65:19]
  wire  soc__T_36; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_32; // @[NutShellSim.scala 65:19]
  wire  soc__T_13; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_31; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_37; // @[NutShellSim.scala 65:19]
  wire  soc__T_26; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_4183; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_4182; // @[NutShellSim.scala 65:19]
  wire  soc__T_33; // @[NutShellSim.scala 65:19]
  wire [63:0] soc__T_4179; // @[NutShellSim.scala 65:19]
  wire  mem_clock; // @[NutShellSim.scala 66:19]
  wire  mem_reset; // @[NutShellSim.scala 66:19]
  wire  mem_io_in_aw_ready; // @[NutShellSim.scala 66:19]
  wire  mem_io_in_aw_valid; // @[NutShellSim.scala 66:19]
  wire [31:0] mem_io_in_aw_bits_addr; // @[NutShellSim.scala 66:19]
  wire  mem_io_in_w_ready; // @[NutShellSim.scala 66:19]
  wire  mem_io_in_w_valid; // @[NutShellSim.scala 66:19]
  wire [63:0] mem_io_in_w_bits_data; // @[NutShellSim.scala 66:19]
  wire  mem_io_in_w_bits_last; // @[NutShellSim.scala 66:19]
  wire  mem_io_in_b_valid; // @[NutShellSim.scala 66:19]
  wire  mem_io_in_ar_ready; // @[NutShellSim.scala 66:19]
  wire  mem_io_in_ar_valid; // @[NutShellSim.scala 66:19]
  wire [31:0] mem_io_in_ar_bits_addr; // @[NutShellSim.scala 66:19]
  wire [7:0] mem_io_in_ar_bits_len; // @[NutShellSim.scala 66:19]
  wire [2:0] mem_io_in_ar_bits_size; // @[NutShellSim.scala 66:19]
  wire [1:0] mem_io_in_ar_bits_burst; // @[NutShellSim.scala 66:19]
  wire  mem_io_in_r_valid; // @[NutShellSim.scala 66:19]
  wire [63:0] mem_io_in_r_bits_data; // @[NutShellSim.scala 66:19]
  wire  mem_io_in_r_bits_last; // @[NutShellSim.scala 66:19]
  wire  memdelay_io_in_aw_ready; // @[NutShellSim.scala 69:24]
  wire  memdelay_io_in_aw_valid; // @[NutShellSim.scala 69:24]
  wire [31:0] memdelay_io_in_aw_bits_addr; // @[NutShellSim.scala 69:24]
  wire [7:0] memdelay_io_in_aw_bits_len; // @[NutShellSim.scala 69:24]
  wire [2:0] memdelay_io_in_aw_bits_size; // @[NutShellSim.scala 69:24]
  wire [1:0] memdelay_io_in_aw_bits_burst; // @[NutShellSim.scala 69:24]
  wire  memdelay_io_in_w_ready; // @[NutShellSim.scala 69:24]
  wire  memdelay_io_in_w_valid; // @[NutShellSim.scala 69:24]
  wire [63:0] memdelay_io_in_w_bits_data; // @[NutShellSim.scala 69:24]
  wire  memdelay_io_in_w_bits_last; // @[NutShellSim.scala 69:24]
  wire  memdelay_io_in_b_valid; // @[NutShellSim.scala 69:24]
  wire  memdelay_io_in_ar_ready; // @[NutShellSim.scala 69:24]
  wire  memdelay_io_in_ar_valid; // @[NutShellSim.scala 69:24]
  wire [31:0] memdelay_io_in_ar_bits_addr; // @[NutShellSim.scala 69:24]
  wire [7:0] memdelay_io_in_ar_bits_len; // @[NutShellSim.scala 69:24]
  wire  memdelay_io_in_r_valid; // @[NutShellSim.scala 69:24]
  wire [63:0] memdelay_io_in_r_bits_data; // @[NutShellSim.scala 69:24]
  wire  memdelay_io_in_r_bits_last; // @[NutShellSim.scala 69:24]
  wire  memdelay_io_out_aw_ready; // @[NutShellSim.scala 69:24]
  wire  memdelay_io_out_aw_valid; // @[NutShellSim.scala 69:24]
  wire [31:0] memdelay_io_out_aw_bits_addr; // @[NutShellSim.scala 69:24]
  wire  memdelay_io_out_w_ready; // @[NutShellSim.scala 69:24]
  wire  memdelay_io_out_w_valid; // @[NutShellSim.scala 69:24]
  wire [63:0] memdelay_io_out_w_bits_data; // @[NutShellSim.scala 69:24]
  wire  memdelay_io_out_w_bits_last; // @[NutShellSim.scala 69:24]
  wire  memdelay_io_out_b_valid; // @[NutShellSim.scala 69:24]
  wire  memdelay_io_out_ar_valid; // @[NutShellSim.scala 69:24]
  wire [31:0] memdelay_io_out_ar_bits_addr; // @[NutShellSim.scala 69:24]
  wire [7:0] memdelay_io_out_ar_bits_len; // @[NutShellSim.scala 69:24]
  wire [2:0] memdelay_io_out_ar_bits_size; // @[NutShellSim.scala 69:24]
  wire [1:0] memdelay_io_out_ar_bits_burst; // @[NutShellSim.scala 69:24]
  wire  memdelay_io_out_r_valid; // @[NutShellSim.scala 69:24]
  wire [63:0] memdelay_io_out_r_bits_data; // @[NutShellSim.scala 69:24]
  wire  memdelay_io_out_r_bits_last; // @[NutShellSim.scala 69:24]
  wire  mmio_clock; // @[NutShellSim.scala 70:20]
  wire  mmio_reset; // @[NutShellSim.scala 70:20]
  wire  mmio_io_rw_req_ready; // @[NutShellSim.scala 70:20]
  wire  mmio_io_rw_req_valid; // @[NutShellSim.scala 70:20]
  wire [31:0] mmio_io_rw_req_bits_addr; // @[NutShellSim.scala 70:20]
  wire [2:0] mmio_io_rw_req_bits_size; // @[NutShellSim.scala 70:20]
  wire [3:0] mmio_io_rw_req_bits_cmd; // @[NutShellSim.scala 70:20]
  wire [7:0] mmio_io_rw_req_bits_wmask; // @[NutShellSim.scala 70:20]
  wire [63:0] mmio_io_rw_req_bits_wdata; // @[NutShellSim.scala 70:20]
  wire  mmio_io_rw_resp_ready; // @[NutShellSim.scala 70:20]
  wire  mmio_io_rw_resp_valid; // @[NutShellSim.scala 70:20]
  wire [63:0] mmio_io_rw_resp_bits_rdata; // @[NutShellSim.scala 70:20]
  wire  mmio_io_difftestCtrl_enable; // @[NutShellSim.scala 70:20]
  wire  mmio_io_meip; // @[NutShellSim.scala 70:20]
  wire  mmio_io_dma_aw_ready; // @[NutShellSim.scala 70:20]
  wire  mmio_io_dma_aw_valid; // @[NutShellSim.scala 70:20]
  wire [31:0] mmio_io_dma_aw_bits_addr; // @[NutShellSim.scala 70:20]
  wire [7:0] mmio_io_dma_aw_bits_len; // @[NutShellSim.scala 70:20]
  wire [2:0] mmio_io_dma_aw_bits_size; // @[NutShellSim.scala 70:20]
  wire  mmio_io_dma_w_ready; // @[NutShellSim.scala 70:20]
  wire  mmio_io_dma_w_valid; // @[NutShellSim.scala 70:20]
  wire [63:0] mmio_io_dma_w_bits_data; // @[NutShellSim.scala 70:20]
  wire [7:0] mmio_io_dma_w_bits_strb; // @[NutShellSim.scala 70:20]
  wire  mmio_io_dma_b_ready; // @[NutShellSim.scala 70:20]
  wire  mmio_io_dma_b_valid; // @[NutShellSim.scala 70:20]
  wire  mmio_io_dma_ar_ready; // @[NutShellSim.scala 70:20]
  wire  mmio_io_dma_ar_valid; // @[NutShellSim.scala 70:20]
  wire [31:0] mmio_io_dma_ar_bits_addr; // @[NutShellSim.scala 70:20]
  wire  mmio_io_dma_r_ready; // @[NutShellSim.scala 70:20]
  wire  mmio_io_dma_r_valid; // @[NutShellSim.scala 70:20]
  wire [63:0] mmio_io_dma_r_bits_data; // @[NutShellSim.scala 70:20]
  wire  mmio__T_13; // @[NutShellSim.scala 70:20]
  wire  _T_1 = io_logCtrl_log_begin <= io_logCtrl_log_end; // @[NutShellSim.scala 105:20]
  wire  _T_3 = _T_1 | reset; // @[NutShellSim.scala 105:9]
  wire  _T_4 = ~_T_3; // @[NutShellSim.scala 105:9]
  reg [63:0] _T_5; // @[GTimer.scala 24:20]
  wire [63:0] _T_7 = _T_5 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_8 = _T_5 >= io_logCtrl_log_begin; // @[NutShellSim.scala 106:35]
  reg [63:0] _T_9; // @[GTimer.scala 24:20]
  wire [63:0] _T_11 = _T_9 + 64'h1; // @[GTimer.scala 25:12]
  wire  _T_12 = _T_9 < io_logCtrl_log_end; // @[NutShellSim.scala 106:62]
  wire  DISPLAY_ENABLE = _T_8 & _T_12; // @[NutShellSim.scala 106:49]
  wire  _T_13 = DISPLAY_ENABLE;
  wire [63:0] difftestThisINST = soc__T_32;
  NutShell soc ( // @[NutShellSim.scala 65:19]
    .clock(soc_clock),
    .reset(soc_reset),
    .io_mem_aw_ready(soc_io_mem_aw_ready),
    .io_mem_aw_valid(soc_io_mem_aw_valid),
    .io_mem_aw_bits_addr(soc_io_mem_aw_bits_addr),
    .io_mem_aw_bits_len(soc_io_mem_aw_bits_len),
    .io_mem_aw_bits_size(soc_io_mem_aw_bits_size),
    .io_mem_aw_bits_burst(soc_io_mem_aw_bits_burst),
    .io_mem_w_ready(soc_io_mem_w_ready),
    .io_mem_w_valid(soc_io_mem_w_valid),
    .io_mem_w_bits_data(soc_io_mem_w_bits_data),
    .io_mem_w_bits_last(soc_io_mem_w_bits_last),
    .io_mem_b_valid(soc_io_mem_b_valid),
    .io_mem_ar_ready(soc_io_mem_ar_ready),
    .io_mem_ar_valid(soc_io_mem_ar_valid),
    .io_mem_ar_bits_addr(soc_io_mem_ar_bits_addr),
    .io_mem_ar_bits_len(soc_io_mem_ar_bits_len),
    .io_mem_r_valid(soc_io_mem_r_valid),
    .io_mem_r_bits_data(soc_io_mem_r_bits_data),
    .io_mem_r_bits_last(soc_io_mem_r_bits_last),
    .io_mmio_req_ready(soc_io_mmio_req_ready),
    .io_mmio_req_valid(soc_io_mmio_req_valid),
    .io_mmio_req_bits_addr(soc_io_mmio_req_bits_addr),
    .io_mmio_req_bits_size(soc_io_mmio_req_bits_size),
    .io_mmio_req_bits_cmd(soc_io_mmio_req_bits_cmd),
    .io_mmio_req_bits_wmask(soc_io_mmio_req_bits_wmask),
    .io_mmio_req_bits_wdata(soc_io_mmio_req_bits_wdata),
    .io_mmio_resp_ready(soc_io_mmio_resp_ready),
    .io_mmio_resp_valid(soc_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(soc_io_mmio_resp_bits_rdata),
    .io_frontend_aw_ready(soc_io_frontend_aw_ready),
    .io_frontend_aw_valid(soc_io_frontend_aw_valid),
    .io_frontend_aw_bits_addr(soc_io_frontend_aw_bits_addr),
    .io_frontend_aw_bits_len(soc_io_frontend_aw_bits_len),
    .io_frontend_aw_bits_size(soc_io_frontend_aw_bits_size),
    .io_frontend_w_ready(soc_io_frontend_w_ready),
    .io_frontend_w_valid(soc_io_frontend_w_valid),
    .io_frontend_w_bits_data(soc_io_frontend_w_bits_data),
    .io_frontend_w_bits_strb(soc_io_frontend_w_bits_strb),
    .io_frontend_b_ready(soc_io_frontend_b_ready),
    .io_frontend_b_valid(soc_io_frontend_b_valid),
    .io_frontend_ar_ready(soc_io_frontend_ar_ready),
    .io_frontend_ar_valid(soc_io_frontend_ar_valid),
    .io_frontend_ar_bits_addr(soc_io_frontend_ar_bits_addr),
    .io_frontend_r_ready(soc_io_frontend_r_ready),
    .io_frontend_r_valid(soc_io_frontend_r_valid),
    .io_frontend_r_bits_data(soc_io_frontend_r_bits_data),
    .io_meip(soc_io_meip),
    ._T_4181(soc__T_4181),
    ._T_4184(soc__T_4184),
    ._T_4185(soc__T_4185),
    .falseWire(soc_falseWire),
    .falseWire_0(soc_falseWire_0),
    ._T_4178(soc__T_4178),
    ._T_284_0(soc__T_284_0),
    ._T_284_1(soc__T_284_1),
    ._T_284_2(soc__T_284_2),
    ._T_284_3(soc__T_284_3),
    ._T_284_4(soc__T_284_4),
    ._T_284_5(soc__T_284_5),
    ._T_284_6(soc__T_284_6),
    ._T_284_7(soc__T_284_7),
    ._T_284_8(soc__T_284_8),
    ._T_284_9(soc__T_284_9),
    ._T_284_10(soc__T_284_10),
    ._T_284_11(soc__T_284_11),
    ._T_284_12(soc__T_284_12),
    ._T_284_13(soc__T_284_13),
    ._T_284_14(soc__T_284_14),
    ._T_284_15(soc__T_284_15),
    ._T_284_16(soc__T_284_16),
    ._T_284_17(soc__T_284_17),
    ._T_284_18(soc__T_284_18),
    ._T_284_19(soc__T_284_19),
    ._T_284_20(soc__T_284_20),
    ._T_284_21(soc__T_284_21),
    ._T_284_22(soc__T_284_22),
    ._T_284_23(soc__T_284_23),
    ._T_284_24(soc__T_284_24),
    ._T_284_25(soc__T_284_25),
    ._T_284_26(soc__T_284_26),
    ._T_284_27(soc__T_284_27),
    ._T_284_28(soc__T_284_28),
    ._T_284_29(soc__T_284_29),
    ._T_284_30(soc__T_284_30),
    ._T_284_31(soc__T_284_31),
    ._T_36(soc__T_36),
    ._T_32(soc__T_32),
    ._T_13(soc__T_13),
    ._T_31(soc__T_31),
    ._T_37(soc__T_37),
    ._T_26(soc__T_26),
    ._T_4183(soc__T_4183),
    ._T_4182(soc__T_4182),
    ._T_33(soc__T_33),
    ._T_4179(soc__T_4179)
  );
  AXI4RAM mem ( // @[NutShellSim.scala 66:19]
    .clock(mem_clock),
    .reset(mem_reset),
    .io_in_aw_ready(mem_io_in_aw_ready),
    .io_in_aw_valid(mem_io_in_aw_valid),
    .io_in_aw_bits_addr(mem_io_in_aw_bits_addr),
    .io_in_w_ready(mem_io_in_w_ready),
    .io_in_w_valid(mem_io_in_w_valid),
    .io_in_w_bits_data(mem_io_in_w_bits_data),
    .io_in_w_bits_last(mem_io_in_w_bits_last),
    .io_in_b_valid(mem_io_in_b_valid),
    .io_in_ar_ready(mem_io_in_ar_ready),
    .io_in_ar_valid(mem_io_in_ar_valid),
    .io_in_ar_bits_addr(mem_io_in_ar_bits_addr),
    .io_in_ar_bits_len(mem_io_in_ar_bits_len),
    .io_in_ar_bits_size(mem_io_in_ar_bits_size),
    .io_in_ar_bits_burst(mem_io_in_ar_bits_burst),
    .io_in_r_valid(mem_io_in_r_valid),
    .io_in_r_bits_data(mem_io_in_r_bits_data),
    .io_in_r_bits_last(mem_io_in_r_bits_last)
  );
  AXI4Delayer memdelay ( // @[NutShellSim.scala 69:24]
    .io_in_aw_ready(memdelay_io_in_aw_ready),
    .io_in_aw_valid(memdelay_io_in_aw_valid),
    .io_in_aw_bits_addr(memdelay_io_in_aw_bits_addr),
    .io_in_aw_bits_len(memdelay_io_in_aw_bits_len),
    .io_in_aw_bits_size(memdelay_io_in_aw_bits_size),
    .io_in_aw_bits_burst(memdelay_io_in_aw_bits_burst),
    .io_in_w_ready(memdelay_io_in_w_ready),
    .io_in_w_valid(memdelay_io_in_w_valid),
    .io_in_w_bits_data(memdelay_io_in_w_bits_data),
    .io_in_w_bits_last(memdelay_io_in_w_bits_last),
    .io_in_b_valid(memdelay_io_in_b_valid),
    .io_in_ar_ready(memdelay_io_in_ar_ready),
    .io_in_ar_valid(memdelay_io_in_ar_valid),
    .io_in_ar_bits_addr(memdelay_io_in_ar_bits_addr),
    .io_in_ar_bits_len(memdelay_io_in_ar_bits_len),
    .io_in_r_valid(memdelay_io_in_r_valid),
    .io_in_r_bits_data(memdelay_io_in_r_bits_data),
    .io_in_r_bits_last(memdelay_io_in_r_bits_last),
    .io_out_aw_ready(memdelay_io_out_aw_ready),
    .io_out_aw_valid(memdelay_io_out_aw_valid),
    .io_out_aw_bits_addr(memdelay_io_out_aw_bits_addr),
    .io_out_w_ready(memdelay_io_out_w_ready),
    .io_out_w_valid(memdelay_io_out_w_valid),
    .io_out_w_bits_data(memdelay_io_out_w_bits_data),
    .io_out_w_bits_last(memdelay_io_out_w_bits_last),
    .io_out_b_valid(memdelay_io_out_b_valid),
    .io_out_ar_valid(memdelay_io_out_ar_valid),
    .io_out_ar_bits_addr(memdelay_io_out_ar_bits_addr),
    .io_out_ar_bits_len(memdelay_io_out_ar_bits_len),
    .io_out_ar_bits_size(memdelay_io_out_ar_bits_size),
    .io_out_ar_bits_burst(memdelay_io_out_ar_bits_burst),
    .io_out_r_valid(memdelay_io_out_r_valid),
    .io_out_r_bits_data(memdelay_io_out_r_bits_data),
    .io_out_r_bits_last(memdelay_io_out_r_bits_last)
  );
  SimMMIO mmio ( // @[NutShellSim.scala 70:20]
    .clock(mmio_clock),
    .reset(mmio_reset),
    .io_rw_req_ready(mmio_io_rw_req_ready),
    .io_rw_req_valid(mmio_io_rw_req_valid),
    .io_rw_req_bits_addr(mmio_io_rw_req_bits_addr),
    .io_rw_req_bits_size(mmio_io_rw_req_bits_size),
    .io_rw_req_bits_cmd(mmio_io_rw_req_bits_cmd),
    .io_rw_req_bits_wmask(mmio_io_rw_req_bits_wmask),
    .io_rw_req_bits_wdata(mmio_io_rw_req_bits_wdata),
    .io_rw_resp_ready(mmio_io_rw_resp_ready),
    .io_rw_resp_valid(mmio_io_rw_resp_valid),
    .io_rw_resp_bits_rdata(mmio_io_rw_resp_bits_rdata),
    .io_difftestCtrl_enable(mmio_io_difftestCtrl_enable),
    .io_meip(mmio_io_meip),
    .io_dma_aw_ready(mmio_io_dma_aw_ready),
    .io_dma_aw_valid(mmio_io_dma_aw_valid),
    .io_dma_aw_bits_addr(mmio_io_dma_aw_bits_addr),
    .io_dma_aw_bits_len(mmio_io_dma_aw_bits_len),
    .io_dma_aw_bits_size(mmio_io_dma_aw_bits_size),
    .io_dma_w_ready(mmio_io_dma_w_ready),
    .io_dma_w_valid(mmio_io_dma_w_valid),
    .io_dma_w_bits_data(mmio_io_dma_w_bits_data),
    .io_dma_w_bits_strb(mmio_io_dma_w_bits_strb),
    .io_dma_b_ready(mmio_io_dma_b_ready),
    .io_dma_b_valid(mmio_io_dma_b_valid),
    .io_dma_ar_ready(mmio_io_dma_ar_ready),
    .io_dma_ar_valid(mmio_io_dma_ar_valid),
    .io_dma_ar_bits_addr(mmio_io_dma_ar_bits_addr),
    .io_dma_r_ready(mmio_io_dma_r_ready),
    .io_dma_r_valid(mmio_io_dma_r_valid),
    .io_dma_r_bits_data(mmio_io_dma_r_bits_data),
    ._T_13(mmio__T_13)
  );
  assign io_difftest_r_0 = soc__T_284_0; // @[NutShellSim.scala 98:15]
  assign io_difftest_r_1 = soc__T_284_1; // @[NutShellSim.scala 98:15]
  assign io_difftest_r_2 = soc__T_284_2; // @[NutShellSim.scala 98:15]
  assign io_difftest_r_3 = soc__T_284_3; // @[NutShellSim.scala 98:15]
  assign io_difftest_r_4 = soc__T_284_4; // @[NutShellSim.scala 98:15]
  assign io_difftest_r_5 = soc__T_284_5; // @[NutShellSim.scala 98:15]
  assign io_difftest_r_6 = soc__T_284_6; // @[NutShellSim.scala 98:15]
  assign io_difftest_r_7 = soc__T_284_7; // @[NutShellSim.scala 98:15]
  assign io_difftest_r_8 = soc__T_284_8; // @[NutShellSim.scala 98:15]
  assign io_difftest_r_9 = soc__T_284_9; // @[NutShellSim.scala 98:15]
  assign io_difftest_r_10 = soc__T_284_10; // @[NutShellSim.scala 98:15]
  assign io_difftest_r_11 = soc__T_284_11; // @[NutShellSim.scala 98:15]
  assign io_difftest_r_12 = soc__T_284_12; // @[NutShellSim.scala 98:15]
  assign io_difftest_r_13 = soc__T_284_13; // @[NutShellSim.scala 98:15]
  assign io_difftest_r_14 = soc__T_284_14; // @[NutShellSim.scala 98:15]
  assign io_difftest_r_15 = soc__T_284_15; // @[NutShellSim.scala 98:15]
  assign io_difftest_r_16 = soc__T_284_16; // @[NutShellSim.scala 98:15]
  assign io_difftest_r_17 = soc__T_284_17; // @[NutShellSim.scala 98:15]
  assign io_difftest_r_18 = soc__T_284_18; // @[NutShellSim.scala 98:15]
  assign io_difftest_r_19 = soc__T_284_19; // @[NutShellSim.scala 98:15]
  assign io_difftest_r_20 = soc__T_284_20; // @[NutShellSim.scala 98:15]
  assign io_difftest_r_21 = soc__T_284_21; // @[NutShellSim.scala 98:15]
  assign io_difftest_r_22 = soc__T_284_22; // @[NutShellSim.scala 98:15]
  assign io_difftest_r_23 = soc__T_284_23; // @[NutShellSim.scala 98:15]
  assign io_difftest_r_24 = soc__T_284_24; // @[NutShellSim.scala 98:15]
  assign io_difftest_r_25 = soc__T_284_25; // @[NutShellSim.scala 98:15]
  assign io_difftest_r_26 = soc__T_284_26; // @[NutShellSim.scala 98:15]
  assign io_difftest_r_27 = soc__T_284_27; // @[NutShellSim.scala 98:15]
  assign io_difftest_r_28 = soc__T_284_28; // @[NutShellSim.scala 98:15]
  assign io_difftest_r_29 = soc__T_284_29; // @[NutShellSim.scala 98:15]
  assign io_difftest_r_30 = soc__T_284_30; // @[NutShellSim.scala 98:15]
  assign io_difftest_r_31 = soc__T_284_31; // @[NutShellSim.scala 98:15]
  assign io_difftest_sr_0 = 64'h0; // @[NutShellSim.scala 98:15]
  assign io_difftest_sr_1 = 64'h0; // @[NutShellSim.scala 98:15]
  assign io_difftest_sr_2 = 64'h0; // @[NutShellSim.scala 98:15]
  assign io_difftest_sr_3 = 64'h0; // @[NutShellSim.scala 98:15]
  assign io_difftest_sr_4 = 64'h0; // @[NutShellSim.scala 98:15]
  assign io_difftest_commit = soc__T_26; // @[NutShellSim.scala 98:15]
  assign io_difftest_isMultiCommit = soc_falseWire; // @[NutShellSim.scala 98:15]
  assign io_difftest_thisPC = soc__T_31; // @[NutShellSim.scala 98:15]
  assign io_difftest_thisINST = difftestThisINST[31:0]; // @[NutShellSim.scala 98:15]
  assign io_difftest_isMMIO = soc__T_33; // @[NutShellSim.scala 98:15]
  assign io_difftest_isRVC = soc__T_36; // @[NutShellSim.scala 98:15]
  assign io_difftest_isRVC2 = soc_falseWire_0; // @[NutShellSim.scala 98:15]
  assign io_difftest_intrNO = soc__T_37; // @[NutShellSim.scala 98:15]
  assign io_difftest_priviledgeMode = soc__T_4178; // @[NutShellSim.scala 98:15]
  assign io_difftest_mstatus = soc__T_4179; // @[NutShellSim.scala 98:15]
  assign io_difftest_sstatus = soc__T_4181; // @[NutShellSim.scala 98:15]
  assign io_difftest_mepc = soc__T_4182; // @[NutShellSim.scala 98:15]
  assign io_difftest_sepc = soc__T_4183; // @[NutShellSim.scala 98:15]
  assign io_difftest_mcause = soc__T_4184; // @[NutShellSim.scala 98:15]
  assign io_difftest_scause = soc__T_4185; // @[NutShellSim.scala 98:15]
  assign io_difftestCtrl_enable = mmio_io_difftestCtrl_enable; // @[NutShellSim.scala 112:19]
  assign soc_clock = clock;
  assign soc_reset = reset;
  assign soc_io_mem_aw_ready = memdelay_io_in_aw_ready; // @[NutShellSim.scala 74:18]
  assign soc_io_mem_w_ready = memdelay_io_in_w_ready; // @[NutShellSim.scala 74:18]
  assign soc_io_mem_b_valid = memdelay_io_in_b_valid; // @[NutShellSim.scala 74:18]
  assign soc_io_mem_ar_ready = memdelay_io_in_ar_ready; // @[NutShellSim.scala 74:18]
  assign soc_io_mem_r_valid = memdelay_io_in_r_valid; // @[NutShellSim.scala 74:18]
  assign soc_io_mem_r_bits_data = memdelay_io_in_r_bits_data; // @[NutShellSim.scala 74:18]
  assign soc_io_mem_r_bits_last = memdelay_io_in_r_bits_last; // @[NutShellSim.scala 74:18]
  assign soc_io_mmio_req_ready = mmio_io_rw_req_ready; // @[NutShellSim.scala 77:14]
  assign soc_io_mmio_resp_valid = mmio_io_rw_resp_valid; // @[NutShellSim.scala 77:14]
  assign soc_io_mmio_resp_bits_rdata = mmio_io_rw_resp_bits_rdata; // @[NutShellSim.scala 77:14]
  assign soc_io_frontend_aw_valid = mmio_io_dma_aw_valid; // @[NutShellSim.scala 72:19]
  assign soc_io_frontend_aw_bits_addr = mmio_io_dma_aw_bits_addr; // @[NutShellSim.scala 72:19]
  assign soc_io_frontend_aw_bits_len = mmio_io_dma_aw_bits_len; // @[NutShellSim.scala 72:19]
  assign soc_io_frontend_aw_bits_size = mmio_io_dma_aw_bits_size; // @[NutShellSim.scala 72:19]
  assign soc_io_frontend_w_valid = mmio_io_dma_w_valid; // @[NutShellSim.scala 72:19]
  assign soc_io_frontend_w_bits_data = mmio_io_dma_w_bits_data; // @[NutShellSim.scala 72:19]
  assign soc_io_frontend_w_bits_strb = mmio_io_dma_w_bits_strb; // @[NutShellSim.scala 72:19]
  assign soc_io_frontend_b_ready = mmio_io_dma_b_ready; // @[NutShellSim.scala 72:19]
  assign soc_io_frontend_ar_valid = mmio_io_dma_ar_valid; // @[NutShellSim.scala 72:19]
  assign soc_io_frontend_ar_bits_addr = mmio_io_dma_ar_bits_addr; // @[NutShellSim.scala 72:19]
  assign soc_io_frontend_r_ready = mmio_io_dma_r_ready; // @[NutShellSim.scala 72:19]
  assign soc_io_meip = mmio_io_meip; // @[NutShellSim.scala 79:15]
  assign soc__T_13 = _T_8 & _T_12;
  assign mem_clock = clock;
  assign mem_reset = reset;
  assign mem_io_in_aw_valid = memdelay_io_out_aw_valid; // @[NutShellSim.scala 75:13]
  assign mem_io_in_aw_bits_addr = memdelay_io_out_aw_bits_addr; // @[NutShellSim.scala 75:13]
  assign mem_io_in_w_valid = memdelay_io_out_w_valid; // @[NutShellSim.scala 75:13]
  assign mem_io_in_w_bits_data = memdelay_io_out_w_bits_data; // @[NutShellSim.scala 75:13]
  assign mem_io_in_w_bits_last = memdelay_io_out_w_bits_last; // @[NutShellSim.scala 75:13]
  assign mem_io_in_ar_valid = memdelay_io_out_ar_valid; // @[NutShellSim.scala 75:13]
  assign mem_io_in_ar_bits_addr = memdelay_io_out_ar_bits_addr; // @[NutShellSim.scala 75:13]
  assign mem_io_in_ar_bits_len = memdelay_io_out_ar_bits_len; // @[NutShellSim.scala 75:13]
  assign mem_io_in_ar_bits_size = memdelay_io_out_ar_bits_size; // @[NutShellSim.scala 75:13]
  assign mem_io_in_ar_bits_burst = memdelay_io_out_ar_bits_burst; // @[NutShellSim.scala 75:13]
  assign memdelay_io_in_aw_valid = soc_io_mem_aw_valid; // @[NutShellSim.scala 74:18]
  assign memdelay_io_in_aw_bits_addr = soc_io_mem_aw_bits_addr; // @[NutShellSim.scala 74:18]
  assign memdelay_io_in_aw_bits_len = soc_io_mem_aw_bits_len; // @[NutShellSim.scala 74:18]
  assign memdelay_io_in_aw_bits_size = soc_io_mem_aw_bits_size; // @[NutShellSim.scala 74:18]
  assign memdelay_io_in_aw_bits_burst = soc_io_mem_aw_bits_burst; // @[NutShellSim.scala 74:18]
  assign memdelay_io_in_w_valid = soc_io_mem_w_valid; // @[NutShellSim.scala 74:18]
  assign memdelay_io_in_w_bits_data = soc_io_mem_w_bits_data; // @[NutShellSim.scala 74:18]
  assign memdelay_io_in_w_bits_last = soc_io_mem_w_bits_last; // @[NutShellSim.scala 74:18]
  assign memdelay_io_in_ar_valid = soc_io_mem_ar_valid; // @[NutShellSim.scala 74:18]
  assign memdelay_io_in_ar_bits_addr = soc_io_mem_ar_bits_addr; // @[NutShellSim.scala 74:18]
  assign memdelay_io_in_ar_bits_len = soc_io_mem_ar_bits_len; // @[NutShellSim.scala 74:18]
  assign memdelay_io_out_aw_ready = mem_io_in_aw_ready; // @[NutShellSim.scala 75:13]
  assign memdelay_io_out_w_ready = mem_io_in_w_ready; // @[NutShellSim.scala 75:13]
  assign memdelay_io_out_b_valid = mem_io_in_b_valid; // @[NutShellSim.scala 75:13]
  assign memdelay_io_out_r_valid = mem_io_in_r_valid; // @[NutShellSim.scala 75:13]
  assign memdelay_io_out_r_bits_data = mem_io_in_r_bits_data; // @[NutShellSim.scala 75:13]
  assign memdelay_io_out_r_bits_last = mem_io_in_r_bits_last; // @[NutShellSim.scala 75:13]
  assign mmio_clock = clock;
  assign mmio_reset = reset;
  assign mmio_io_rw_req_valid = soc_io_mmio_req_valid; // @[NutShellSim.scala 77:14]
  assign mmio_io_rw_req_bits_addr = soc_io_mmio_req_bits_addr; // @[NutShellSim.scala 77:14]
  assign mmio_io_rw_req_bits_size = soc_io_mmio_req_bits_size; // @[NutShellSim.scala 77:14]
  assign mmio_io_rw_req_bits_cmd = soc_io_mmio_req_bits_cmd; // @[NutShellSim.scala 77:14]
  assign mmio_io_rw_req_bits_wmask = soc_io_mmio_req_bits_wmask; // @[NutShellSim.scala 77:14]
  assign mmio_io_rw_req_bits_wdata = soc_io_mmio_req_bits_wdata; // @[NutShellSim.scala 77:14]
  assign mmio_io_rw_resp_ready = soc_io_mmio_resp_ready; // @[NutShellSim.scala 77:14]
  assign mmio_io_dma_aw_ready = soc_io_frontend_aw_ready; // @[NutShellSim.scala 72:19]
  assign mmio_io_dma_w_ready = soc_io_frontend_w_ready; // @[NutShellSim.scala 72:19]
  assign mmio_io_dma_b_valid = soc_io_frontend_b_valid; // @[NutShellSim.scala 72:19]
  assign mmio_io_dma_ar_ready = soc_io_frontend_ar_ready; // @[NutShellSim.scala 72:19]
  assign mmio_io_dma_r_valid = soc_io_frontend_r_valid; // @[NutShellSim.scala 72:19]
  assign mmio_io_dma_r_bits_data = soc_io_frontend_r_bits_data; // @[NutShellSim.scala 72:19]
  assign mmio__T_13 = _T_8 & _T_12;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  _T_5 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  _T_9 = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_5 <= 64'h0;
    end else begin
      _T_5 <= _T_7;
    end
    if (reset) begin
      _T_9 <= 64'h0;
    end else begin
      _T_9 <= _T_11;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4) begin
          $fwrite(32'h80000002,"Assertion failed\n    at NutShellSim.scala:105 assert(log_begin <= log_end)\n"); // @[NutShellSim.scala 105:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_4) begin
          $fatal; // @[NutShellSim.scala 105:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
